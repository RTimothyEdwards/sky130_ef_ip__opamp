magic
tech sky130A
magscale 1 2
timestamp 1652924542
<< pwell >>
rect -3359 -776 3359 776
<< mvnmos >>
rect -3131 318 -3031 518
rect -2973 318 -2873 518
rect -2815 318 -2715 518
rect -2657 318 -2557 518
rect -2499 318 -2399 518
rect -2341 318 -2241 518
rect -2183 318 -2083 518
rect -2025 318 -1925 518
rect -1867 318 -1767 518
rect -1709 318 -1609 518
rect -1551 318 -1451 518
rect -1393 318 -1293 518
rect -1235 318 -1135 518
rect -1077 318 -977 518
rect -919 318 -819 518
rect -761 318 -661 518
rect -603 318 -503 518
rect -445 318 -345 518
rect -287 318 -187 518
rect -129 318 -29 518
rect 29 318 129 518
rect 187 318 287 518
rect 345 318 445 518
rect 503 318 603 518
rect 661 318 761 518
rect 819 318 919 518
rect 977 318 1077 518
rect 1135 318 1235 518
rect 1293 318 1393 518
rect 1451 318 1551 518
rect 1609 318 1709 518
rect 1767 318 1867 518
rect 1925 318 2025 518
rect 2083 318 2183 518
rect 2241 318 2341 518
rect 2399 318 2499 518
rect 2557 318 2657 518
rect 2715 318 2815 518
rect 2873 318 2973 518
rect 3031 318 3131 518
rect -3131 -100 -3031 100
rect -2973 -100 -2873 100
rect -2815 -100 -2715 100
rect -2657 -100 -2557 100
rect -2499 -100 -2399 100
rect -2341 -100 -2241 100
rect -2183 -100 -2083 100
rect -2025 -100 -1925 100
rect -1867 -100 -1767 100
rect -1709 -100 -1609 100
rect -1551 -100 -1451 100
rect -1393 -100 -1293 100
rect -1235 -100 -1135 100
rect -1077 -100 -977 100
rect -919 -100 -819 100
rect -761 -100 -661 100
rect -603 -100 -503 100
rect -445 -100 -345 100
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
rect 345 -100 445 100
rect 503 -100 603 100
rect 661 -100 761 100
rect 819 -100 919 100
rect 977 -100 1077 100
rect 1135 -100 1235 100
rect 1293 -100 1393 100
rect 1451 -100 1551 100
rect 1609 -100 1709 100
rect 1767 -100 1867 100
rect 1925 -100 2025 100
rect 2083 -100 2183 100
rect 2241 -100 2341 100
rect 2399 -100 2499 100
rect 2557 -100 2657 100
rect 2715 -100 2815 100
rect 2873 -100 2973 100
rect 3031 -100 3131 100
rect -3131 -518 -3031 -318
rect -2973 -518 -2873 -318
rect -2815 -518 -2715 -318
rect -2657 -518 -2557 -318
rect -2499 -518 -2399 -318
rect -2341 -518 -2241 -318
rect -2183 -518 -2083 -318
rect -2025 -518 -1925 -318
rect -1867 -518 -1767 -318
rect -1709 -518 -1609 -318
rect -1551 -518 -1451 -318
rect -1393 -518 -1293 -318
rect -1235 -518 -1135 -318
rect -1077 -518 -977 -318
rect -919 -518 -819 -318
rect -761 -518 -661 -318
rect -603 -518 -503 -318
rect -445 -518 -345 -318
rect -287 -518 -187 -318
rect -129 -518 -29 -318
rect 29 -518 129 -318
rect 187 -518 287 -318
rect 345 -518 445 -318
rect 503 -518 603 -318
rect 661 -518 761 -318
rect 819 -518 919 -318
rect 977 -518 1077 -318
rect 1135 -518 1235 -318
rect 1293 -518 1393 -318
rect 1451 -518 1551 -318
rect 1609 -518 1709 -318
rect 1767 -518 1867 -318
rect 1925 -518 2025 -318
rect 2083 -518 2183 -318
rect 2241 -518 2341 -318
rect 2399 -518 2499 -318
rect 2557 -518 2657 -318
rect 2715 -518 2815 -318
rect 2873 -518 2973 -318
rect 3031 -518 3131 -318
<< mvndiff >>
rect -3189 506 -3131 518
rect -3189 330 -3177 506
rect -3143 330 -3131 506
rect -3189 318 -3131 330
rect -3031 506 -2973 518
rect -3031 330 -3019 506
rect -2985 330 -2973 506
rect -3031 318 -2973 330
rect -2873 506 -2815 518
rect -2873 330 -2861 506
rect -2827 330 -2815 506
rect -2873 318 -2815 330
rect -2715 506 -2657 518
rect -2715 330 -2703 506
rect -2669 330 -2657 506
rect -2715 318 -2657 330
rect -2557 506 -2499 518
rect -2557 330 -2545 506
rect -2511 330 -2499 506
rect -2557 318 -2499 330
rect -2399 506 -2341 518
rect -2399 330 -2387 506
rect -2353 330 -2341 506
rect -2399 318 -2341 330
rect -2241 506 -2183 518
rect -2241 330 -2229 506
rect -2195 330 -2183 506
rect -2241 318 -2183 330
rect -2083 506 -2025 518
rect -2083 330 -2071 506
rect -2037 330 -2025 506
rect -2083 318 -2025 330
rect -1925 506 -1867 518
rect -1925 330 -1913 506
rect -1879 330 -1867 506
rect -1925 318 -1867 330
rect -1767 506 -1709 518
rect -1767 330 -1755 506
rect -1721 330 -1709 506
rect -1767 318 -1709 330
rect -1609 506 -1551 518
rect -1609 330 -1597 506
rect -1563 330 -1551 506
rect -1609 318 -1551 330
rect -1451 506 -1393 518
rect -1451 330 -1439 506
rect -1405 330 -1393 506
rect -1451 318 -1393 330
rect -1293 506 -1235 518
rect -1293 330 -1281 506
rect -1247 330 -1235 506
rect -1293 318 -1235 330
rect -1135 506 -1077 518
rect -1135 330 -1123 506
rect -1089 330 -1077 506
rect -1135 318 -1077 330
rect -977 506 -919 518
rect -977 330 -965 506
rect -931 330 -919 506
rect -977 318 -919 330
rect -819 506 -761 518
rect -819 330 -807 506
rect -773 330 -761 506
rect -819 318 -761 330
rect -661 506 -603 518
rect -661 330 -649 506
rect -615 330 -603 506
rect -661 318 -603 330
rect -503 506 -445 518
rect -503 330 -491 506
rect -457 330 -445 506
rect -503 318 -445 330
rect -345 506 -287 518
rect -345 330 -333 506
rect -299 330 -287 506
rect -345 318 -287 330
rect -187 506 -129 518
rect -187 330 -175 506
rect -141 330 -129 506
rect -187 318 -129 330
rect -29 506 29 518
rect -29 330 -17 506
rect 17 330 29 506
rect -29 318 29 330
rect 129 506 187 518
rect 129 330 141 506
rect 175 330 187 506
rect 129 318 187 330
rect 287 506 345 518
rect 287 330 299 506
rect 333 330 345 506
rect 287 318 345 330
rect 445 506 503 518
rect 445 330 457 506
rect 491 330 503 506
rect 445 318 503 330
rect 603 506 661 518
rect 603 330 615 506
rect 649 330 661 506
rect 603 318 661 330
rect 761 506 819 518
rect 761 330 773 506
rect 807 330 819 506
rect 761 318 819 330
rect 919 506 977 518
rect 919 330 931 506
rect 965 330 977 506
rect 919 318 977 330
rect 1077 506 1135 518
rect 1077 330 1089 506
rect 1123 330 1135 506
rect 1077 318 1135 330
rect 1235 506 1293 518
rect 1235 330 1247 506
rect 1281 330 1293 506
rect 1235 318 1293 330
rect 1393 506 1451 518
rect 1393 330 1405 506
rect 1439 330 1451 506
rect 1393 318 1451 330
rect 1551 506 1609 518
rect 1551 330 1563 506
rect 1597 330 1609 506
rect 1551 318 1609 330
rect 1709 506 1767 518
rect 1709 330 1721 506
rect 1755 330 1767 506
rect 1709 318 1767 330
rect 1867 506 1925 518
rect 1867 330 1879 506
rect 1913 330 1925 506
rect 1867 318 1925 330
rect 2025 506 2083 518
rect 2025 330 2037 506
rect 2071 330 2083 506
rect 2025 318 2083 330
rect 2183 506 2241 518
rect 2183 330 2195 506
rect 2229 330 2241 506
rect 2183 318 2241 330
rect 2341 506 2399 518
rect 2341 330 2353 506
rect 2387 330 2399 506
rect 2341 318 2399 330
rect 2499 506 2557 518
rect 2499 330 2511 506
rect 2545 330 2557 506
rect 2499 318 2557 330
rect 2657 506 2715 518
rect 2657 330 2669 506
rect 2703 330 2715 506
rect 2657 318 2715 330
rect 2815 506 2873 518
rect 2815 330 2827 506
rect 2861 330 2873 506
rect 2815 318 2873 330
rect 2973 506 3031 518
rect 2973 330 2985 506
rect 3019 330 3031 506
rect 2973 318 3031 330
rect 3131 506 3189 518
rect 3131 330 3143 506
rect 3177 330 3189 506
rect 3131 318 3189 330
rect -3189 88 -3131 100
rect -3189 -88 -3177 88
rect -3143 -88 -3131 88
rect -3189 -100 -3131 -88
rect -3031 88 -2973 100
rect -3031 -88 -3019 88
rect -2985 -88 -2973 88
rect -3031 -100 -2973 -88
rect -2873 88 -2815 100
rect -2873 -88 -2861 88
rect -2827 -88 -2815 88
rect -2873 -100 -2815 -88
rect -2715 88 -2657 100
rect -2715 -88 -2703 88
rect -2669 -88 -2657 88
rect -2715 -100 -2657 -88
rect -2557 88 -2499 100
rect -2557 -88 -2545 88
rect -2511 -88 -2499 88
rect -2557 -100 -2499 -88
rect -2399 88 -2341 100
rect -2399 -88 -2387 88
rect -2353 -88 -2341 88
rect -2399 -100 -2341 -88
rect -2241 88 -2183 100
rect -2241 -88 -2229 88
rect -2195 -88 -2183 88
rect -2241 -100 -2183 -88
rect -2083 88 -2025 100
rect -2083 -88 -2071 88
rect -2037 -88 -2025 88
rect -2083 -100 -2025 -88
rect -1925 88 -1867 100
rect -1925 -88 -1913 88
rect -1879 -88 -1867 88
rect -1925 -100 -1867 -88
rect -1767 88 -1709 100
rect -1767 -88 -1755 88
rect -1721 -88 -1709 88
rect -1767 -100 -1709 -88
rect -1609 88 -1551 100
rect -1609 -88 -1597 88
rect -1563 -88 -1551 88
rect -1609 -100 -1551 -88
rect -1451 88 -1393 100
rect -1451 -88 -1439 88
rect -1405 -88 -1393 88
rect -1451 -100 -1393 -88
rect -1293 88 -1235 100
rect -1293 -88 -1281 88
rect -1247 -88 -1235 88
rect -1293 -100 -1235 -88
rect -1135 88 -1077 100
rect -1135 -88 -1123 88
rect -1089 -88 -1077 88
rect -1135 -100 -1077 -88
rect -977 88 -919 100
rect -977 -88 -965 88
rect -931 -88 -919 88
rect -977 -100 -919 -88
rect -819 88 -761 100
rect -819 -88 -807 88
rect -773 -88 -761 88
rect -819 -100 -761 -88
rect -661 88 -603 100
rect -661 -88 -649 88
rect -615 -88 -603 88
rect -661 -100 -603 -88
rect -503 88 -445 100
rect -503 -88 -491 88
rect -457 -88 -445 88
rect -503 -100 -445 -88
rect -345 88 -287 100
rect -345 -88 -333 88
rect -299 -88 -287 88
rect -345 -100 -287 -88
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
rect 287 88 345 100
rect 287 -88 299 88
rect 333 -88 345 88
rect 287 -100 345 -88
rect 445 88 503 100
rect 445 -88 457 88
rect 491 -88 503 88
rect 445 -100 503 -88
rect 603 88 661 100
rect 603 -88 615 88
rect 649 -88 661 88
rect 603 -100 661 -88
rect 761 88 819 100
rect 761 -88 773 88
rect 807 -88 819 88
rect 761 -100 819 -88
rect 919 88 977 100
rect 919 -88 931 88
rect 965 -88 977 88
rect 919 -100 977 -88
rect 1077 88 1135 100
rect 1077 -88 1089 88
rect 1123 -88 1135 88
rect 1077 -100 1135 -88
rect 1235 88 1293 100
rect 1235 -88 1247 88
rect 1281 -88 1293 88
rect 1235 -100 1293 -88
rect 1393 88 1451 100
rect 1393 -88 1405 88
rect 1439 -88 1451 88
rect 1393 -100 1451 -88
rect 1551 88 1609 100
rect 1551 -88 1563 88
rect 1597 -88 1609 88
rect 1551 -100 1609 -88
rect 1709 88 1767 100
rect 1709 -88 1721 88
rect 1755 -88 1767 88
rect 1709 -100 1767 -88
rect 1867 88 1925 100
rect 1867 -88 1879 88
rect 1913 -88 1925 88
rect 1867 -100 1925 -88
rect 2025 88 2083 100
rect 2025 -88 2037 88
rect 2071 -88 2083 88
rect 2025 -100 2083 -88
rect 2183 88 2241 100
rect 2183 -88 2195 88
rect 2229 -88 2241 88
rect 2183 -100 2241 -88
rect 2341 88 2399 100
rect 2341 -88 2353 88
rect 2387 -88 2399 88
rect 2341 -100 2399 -88
rect 2499 88 2557 100
rect 2499 -88 2511 88
rect 2545 -88 2557 88
rect 2499 -100 2557 -88
rect 2657 88 2715 100
rect 2657 -88 2669 88
rect 2703 -88 2715 88
rect 2657 -100 2715 -88
rect 2815 88 2873 100
rect 2815 -88 2827 88
rect 2861 -88 2873 88
rect 2815 -100 2873 -88
rect 2973 88 3031 100
rect 2973 -88 2985 88
rect 3019 -88 3031 88
rect 2973 -100 3031 -88
rect 3131 88 3189 100
rect 3131 -88 3143 88
rect 3177 -88 3189 88
rect 3131 -100 3189 -88
rect -3189 -330 -3131 -318
rect -3189 -506 -3177 -330
rect -3143 -506 -3131 -330
rect -3189 -518 -3131 -506
rect -3031 -330 -2973 -318
rect -3031 -506 -3019 -330
rect -2985 -506 -2973 -330
rect -3031 -518 -2973 -506
rect -2873 -330 -2815 -318
rect -2873 -506 -2861 -330
rect -2827 -506 -2815 -330
rect -2873 -518 -2815 -506
rect -2715 -330 -2657 -318
rect -2715 -506 -2703 -330
rect -2669 -506 -2657 -330
rect -2715 -518 -2657 -506
rect -2557 -330 -2499 -318
rect -2557 -506 -2545 -330
rect -2511 -506 -2499 -330
rect -2557 -518 -2499 -506
rect -2399 -330 -2341 -318
rect -2399 -506 -2387 -330
rect -2353 -506 -2341 -330
rect -2399 -518 -2341 -506
rect -2241 -330 -2183 -318
rect -2241 -506 -2229 -330
rect -2195 -506 -2183 -330
rect -2241 -518 -2183 -506
rect -2083 -330 -2025 -318
rect -2083 -506 -2071 -330
rect -2037 -506 -2025 -330
rect -2083 -518 -2025 -506
rect -1925 -330 -1867 -318
rect -1925 -506 -1913 -330
rect -1879 -506 -1867 -330
rect -1925 -518 -1867 -506
rect -1767 -330 -1709 -318
rect -1767 -506 -1755 -330
rect -1721 -506 -1709 -330
rect -1767 -518 -1709 -506
rect -1609 -330 -1551 -318
rect -1609 -506 -1597 -330
rect -1563 -506 -1551 -330
rect -1609 -518 -1551 -506
rect -1451 -330 -1393 -318
rect -1451 -506 -1439 -330
rect -1405 -506 -1393 -330
rect -1451 -518 -1393 -506
rect -1293 -330 -1235 -318
rect -1293 -506 -1281 -330
rect -1247 -506 -1235 -330
rect -1293 -518 -1235 -506
rect -1135 -330 -1077 -318
rect -1135 -506 -1123 -330
rect -1089 -506 -1077 -330
rect -1135 -518 -1077 -506
rect -977 -330 -919 -318
rect -977 -506 -965 -330
rect -931 -506 -919 -330
rect -977 -518 -919 -506
rect -819 -330 -761 -318
rect -819 -506 -807 -330
rect -773 -506 -761 -330
rect -819 -518 -761 -506
rect -661 -330 -603 -318
rect -661 -506 -649 -330
rect -615 -506 -603 -330
rect -661 -518 -603 -506
rect -503 -330 -445 -318
rect -503 -506 -491 -330
rect -457 -506 -445 -330
rect -503 -518 -445 -506
rect -345 -330 -287 -318
rect -345 -506 -333 -330
rect -299 -506 -287 -330
rect -345 -518 -287 -506
rect -187 -330 -129 -318
rect -187 -506 -175 -330
rect -141 -506 -129 -330
rect -187 -518 -129 -506
rect -29 -330 29 -318
rect -29 -506 -17 -330
rect 17 -506 29 -330
rect -29 -518 29 -506
rect 129 -330 187 -318
rect 129 -506 141 -330
rect 175 -506 187 -330
rect 129 -518 187 -506
rect 287 -330 345 -318
rect 287 -506 299 -330
rect 333 -506 345 -330
rect 287 -518 345 -506
rect 445 -330 503 -318
rect 445 -506 457 -330
rect 491 -506 503 -330
rect 445 -518 503 -506
rect 603 -330 661 -318
rect 603 -506 615 -330
rect 649 -506 661 -330
rect 603 -518 661 -506
rect 761 -330 819 -318
rect 761 -506 773 -330
rect 807 -506 819 -330
rect 761 -518 819 -506
rect 919 -330 977 -318
rect 919 -506 931 -330
rect 965 -506 977 -330
rect 919 -518 977 -506
rect 1077 -330 1135 -318
rect 1077 -506 1089 -330
rect 1123 -506 1135 -330
rect 1077 -518 1135 -506
rect 1235 -330 1293 -318
rect 1235 -506 1247 -330
rect 1281 -506 1293 -330
rect 1235 -518 1293 -506
rect 1393 -330 1451 -318
rect 1393 -506 1405 -330
rect 1439 -506 1451 -330
rect 1393 -518 1451 -506
rect 1551 -330 1609 -318
rect 1551 -506 1563 -330
rect 1597 -506 1609 -330
rect 1551 -518 1609 -506
rect 1709 -330 1767 -318
rect 1709 -506 1721 -330
rect 1755 -506 1767 -330
rect 1709 -518 1767 -506
rect 1867 -330 1925 -318
rect 1867 -506 1879 -330
rect 1913 -506 1925 -330
rect 1867 -518 1925 -506
rect 2025 -330 2083 -318
rect 2025 -506 2037 -330
rect 2071 -506 2083 -330
rect 2025 -518 2083 -506
rect 2183 -330 2241 -318
rect 2183 -506 2195 -330
rect 2229 -506 2241 -330
rect 2183 -518 2241 -506
rect 2341 -330 2399 -318
rect 2341 -506 2353 -330
rect 2387 -506 2399 -330
rect 2341 -518 2399 -506
rect 2499 -330 2557 -318
rect 2499 -506 2511 -330
rect 2545 -506 2557 -330
rect 2499 -518 2557 -506
rect 2657 -330 2715 -318
rect 2657 -506 2669 -330
rect 2703 -506 2715 -330
rect 2657 -518 2715 -506
rect 2815 -330 2873 -318
rect 2815 -506 2827 -330
rect 2861 -506 2873 -330
rect 2815 -518 2873 -506
rect 2973 -330 3031 -318
rect 2973 -506 2985 -330
rect 3019 -506 3031 -330
rect 2973 -518 3031 -506
rect 3131 -330 3189 -318
rect 3131 -506 3143 -330
rect 3177 -506 3189 -330
rect 3131 -518 3189 -506
<< mvndiffc >>
rect -3177 330 -3143 506
rect -3019 330 -2985 506
rect -2861 330 -2827 506
rect -2703 330 -2669 506
rect -2545 330 -2511 506
rect -2387 330 -2353 506
rect -2229 330 -2195 506
rect -2071 330 -2037 506
rect -1913 330 -1879 506
rect -1755 330 -1721 506
rect -1597 330 -1563 506
rect -1439 330 -1405 506
rect -1281 330 -1247 506
rect -1123 330 -1089 506
rect -965 330 -931 506
rect -807 330 -773 506
rect -649 330 -615 506
rect -491 330 -457 506
rect -333 330 -299 506
rect -175 330 -141 506
rect -17 330 17 506
rect 141 330 175 506
rect 299 330 333 506
rect 457 330 491 506
rect 615 330 649 506
rect 773 330 807 506
rect 931 330 965 506
rect 1089 330 1123 506
rect 1247 330 1281 506
rect 1405 330 1439 506
rect 1563 330 1597 506
rect 1721 330 1755 506
rect 1879 330 1913 506
rect 2037 330 2071 506
rect 2195 330 2229 506
rect 2353 330 2387 506
rect 2511 330 2545 506
rect 2669 330 2703 506
rect 2827 330 2861 506
rect 2985 330 3019 506
rect 3143 330 3177 506
rect -3177 -88 -3143 88
rect -3019 -88 -2985 88
rect -2861 -88 -2827 88
rect -2703 -88 -2669 88
rect -2545 -88 -2511 88
rect -2387 -88 -2353 88
rect -2229 -88 -2195 88
rect -2071 -88 -2037 88
rect -1913 -88 -1879 88
rect -1755 -88 -1721 88
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
rect 1721 -88 1755 88
rect 1879 -88 1913 88
rect 2037 -88 2071 88
rect 2195 -88 2229 88
rect 2353 -88 2387 88
rect 2511 -88 2545 88
rect 2669 -88 2703 88
rect 2827 -88 2861 88
rect 2985 -88 3019 88
rect 3143 -88 3177 88
rect -3177 -506 -3143 -330
rect -3019 -506 -2985 -330
rect -2861 -506 -2827 -330
rect -2703 -506 -2669 -330
rect -2545 -506 -2511 -330
rect -2387 -506 -2353 -330
rect -2229 -506 -2195 -330
rect -2071 -506 -2037 -330
rect -1913 -506 -1879 -330
rect -1755 -506 -1721 -330
rect -1597 -506 -1563 -330
rect -1439 -506 -1405 -330
rect -1281 -506 -1247 -330
rect -1123 -506 -1089 -330
rect -965 -506 -931 -330
rect -807 -506 -773 -330
rect -649 -506 -615 -330
rect -491 -506 -457 -330
rect -333 -506 -299 -330
rect -175 -506 -141 -330
rect -17 -506 17 -330
rect 141 -506 175 -330
rect 299 -506 333 -330
rect 457 -506 491 -330
rect 615 -506 649 -330
rect 773 -506 807 -330
rect 931 -506 965 -330
rect 1089 -506 1123 -330
rect 1247 -506 1281 -330
rect 1405 -506 1439 -330
rect 1563 -506 1597 -330
rect 1721 -506 1755 -330
rect 1879 -506 1913 -330
rect 2037 -506 2071 -330
rect 2195 -506 2229 -330
rect 2353 -506 2387 -330
rect 2511 -506 2545 -330
rect 2669 -506 2703 -330
rect 2827 -506 2861 -330
rect 2985 -506 3019 -330
rect 3143 -506 3177 -330
<< mvpsubdiff >>
rect -3323 728 3323 740
rect -3323 694 -3215 728
rect 3215 694 3323 728
rect -3323 682 3323 694
rect -3323 632 -3265 682
rect -3323 -632 -3311 632
rect -3277 -632 -3265 632
rect 3265 632 3323 682
rect -3323 -682 -3265 -632
rect 3265 -632 3277 632
rect 3311 -632 3323 632
rect 3265 -682 3323 -632
rect -3323 -694 3323 -682
rect -3323 -728 -3215 -694
rect 3215 -728 3323 -694
rect -3323 -740 3323 -728
<< mvpsubdiffcont >>
rect -3215 694 3215 728
rect -3311 -632 -3277 632
rect 3277 -632 3311 632
rect -3215 -728 3215 -694
<< poly >>
rect -3131 590 -3031 606
rect -3131 556 -3115 590
rect -3047 556 -3031 590
rect -3131 518 -3031 556
rect -2973 590 -2873 606
rect -2973 556 -2957 590
rect -2889 556 -2873 590
rect -2973 518 -2873 556
rect -2815 590 -2715 606
rect -2815 556 -2799 590
rect -2731 556 -2715 590
rect -2815 518 -2715 556
rect -2657 590 -2557 606
rect -2657 556 -2641 590
rect -2573 556 -2557 590
rect -2657 518 -2557 556
rect -2499 590 -2399 606
rect -2499 556 -2483 590
rect -2415 556 -2399 590
rect -2499 518 -2399 556
rect -2341 590 -2241 606
rect -2341 556 -2325 590
rect -2257 556 -2241 590
rect -2341 518 -2241 556
rect -2183 590 -2083 606
rect -2183 556 -2167 590
rect -2099 556 -2083 590
rect -2183 518 -2083 556
rect -2025 590 -1925 606
rect -2025 556 -2009 590
rect -1941 556 -1925 590
rect -2025 518 -1925 556
rect -1867 590 -1767 606
rect -1867 556 -1851 590
rect -1783 556 -1767 590
rect -1867 518 -1767 556
rect -1709 590 -1609 606
rect -1709 556 -1693 590
rect -1625 556 -1609 590
rect -1709 518 -1609 556
rect -1551 590 -1451 606
rect -1551 556 -1535 590
rect -1467 556 -1451 590
rect -1551 518 -1451 556
rect -1393 590 -1293 606
rect -1393 556 -1377 590
rect -1309 556 -1293 590
rect -1393 518 -1293 556
rect -1235 590 -1135 606
rect -1235 556 -1219 590
rect -1151 556 -1135 590
rect -1235 518 -1135 556
rect -1077 590 -977 606
rect -1077 556 -1061 590
rect -993 556 -977 590
rect -1077 518 -977 556
rect -919 590 -819 606
rect -919 556 -903 590
rect -835 556 -819 590
rect -919 518 -819 556
rect -761 590 -661 606
rect -761 556 -745 590
rect -677 556 -661 590
rect -761 518 -661 556
rect -603 590 -503 606
rect -603 556 -587 590
rect -519 556 -503 590
rect -603 518 -503 556
rect -445 590 -345 606
rect -445 556 -429 590
rect -361 556 -345 590
rect -445 518 -345 556
rect -287 590 -187 606
rect -287 556 -271 590
rect -203 556 -187 590
rect -287 518 -187 556
rect -129 590 -29 606
rect -129 556 -113 590
rect -45 556 -29 590
rect -129 518 -29 556
rect 29 590 129 606
rect 29 556 45 590
rect 113 556 129 590
rect 29 518 129 556
rect 187 590 287 606
rect 187 556 203 590
rect 271 556 287 590
rect 187 518 287 556
rect 345 590 445 606
rect 345 556 361 590
rect 429 556 445 590
rect 345 518 445 556
rect 503 590 603 606
rect 503 556 519 590
rect 587 556 603 590
rect 503 518 603 556
rect 661 590 761 606
rect 661 556 677 590
rect 745 556 761 590
rect 661 518 761 556
rect 819 590 919 606
rect 819 556 835 590
rect 903 556 919 590
rect 819 518 919 556
rect 977 590 1077 606
rect 977 556 993 590
rect 1061 556 1077 590
rect 977 518 1077 556
rect 1135 590 1235 606
rect 1135 556 1151 590
rect 1219 556 1235 590
rect 1135 518 1235 556
rect 1293 590 1393 606
rect 1293 556 1309 590
rect 1377 556 1393 590
rect 1293 518 1393 556
rect 1451 590 1551 606
rect 1451 556 1467 590
rect 1535 556 1551 590
rect 1451 518 1551 556
rect 1609 590 1709 606
rect 1609 556 1625 590
rect 1693 556 1709 590
rect 1609 518 1709 556
rect 1767 590 1867 606
rect 1767 556 1783 590
rect 1851 556 1867 590
rect 1767 518 1867 556
rect 1925 590 2025 606
rect 1925 556 1941 590
rect 2009 556 2025 590
rect 1925 518 2025 556
rect 2083 590 2183 606
rect 2083 556 2099 590
rect 2167 556 2183 590
rect 2083 518 2183 556
rect 2241 590 2341 606
rect 2241 556 2257 590
rect 2325 556 2341 590
rect 2241 518 2341 556
rect 2399 590 2499 606
rect 2399 556 2415 590
rect 2483 556 2499 590
rect 2399 518 2499 556
rect 2557 590 2657 606
rect 2557 556 2573 590
rect 2641 556 2657 590
rect 2557 518 2657 556
rect 2715 590 2815 606
rect 2715 556 2731 590
rect 2799 556 2815 590
rect 2715 518 2815 556
rect 2873 590 2973 606
rect 2873 556 2889 590
rect 2957 556 2973 590
rect 2873 518 2973 556
rect 3031 590 3131 606
rect 3031 556 3047 590
rect 3115 556 3131 590
rect 3031 518 3131 556
rect -3131 280 -3031 318
rect -3131 246 -3115 280
rect -3047 246 -3031 280
rect -3131 230 -3031 246
rect -2973 280 -2873 318
rect -2973 246 -2957 280
rect -2889 246 -2873 280
rect -2973 230 -2873 246
rect -2815 280 -2715 318
rect -2815 246 -2799 280
rect -2731 246 -2715 280
rect -2815 230 -2715 246
rect -2657 280 -2557 318
rect -2657 246 -2641 280
rect -2573 246 -2557 280
rect -2657 230 -2557 246
rect -2499 280 -2399 318
rect -2499 246 -2483 280
rect -2415 246 -2399 280
rect -2499 230 -2399 246
rect -2341 280 -2241 318
rect -2341 246 -2325 280
rect -2257 246 -2241 280
rect -2341 230 -2241 246
rect -2183 280 -2083 318
rect -2183 246 -2167 280
rect -2099 246 -2083 280
rect -2183 230 -2083 246
rect -2025 280 -1925 318
rect -2025 246 -2009 280
rect -1941 246 -1925 280
rect -2025 230 -1925 246
rect -1867 280 -1767 318
rect -1867 246 -1851 280
rect -1783 246 -1767 280
rect -1867 230 -1767 246
rect -1709 280 -1609 318
rect -1709 246 -1693 280
rect -1625 246 -1609 280
rect -1709 230 -1609 246
rect -1551 280 -1451 318
rect -1551 246 -1535 280
rect -1467 246 -1451 280
rect -1551 230 -1451 246
rect -1393 280 -1293 318
rect -1393 246 -1377 280
rect -1309 246 -1293 280
rect -1393 230 -1293 246
rect -1235 280 -1135 318
rect -1235 246 -1219 280
rect -1151 246 -1135 280
rect -1235 230 -1135 246
rect -1077 280 -977 318
rect -1077 246 -1061 280
rect -993 246 -977 280
rect -1077 230 -977 246
rect -919 280 -819 318
rect -919 246 -903 280
rect -835 246 -819 280
rect -919 230 -819 246
rect -761 280 -661 318
rect -761 246 -745 280
rect -677 246 -661 280
rect -761 230 -661 246
rect -603 280 -503 318
rect -603 246 -587 280
rect -519 246 -503 280
rect -603 230 -503 246
rect -445 280 -345 318
rect -445 246 -429 280
rect -361 246 -345 280
rect -445 230 -345 246
rect -287 280 -187 318
rect -287 246 -271 280
rect -203 246 -187 280
rect -287 230 -187 246
rect -129 280 -29 318
rect -129 246 -113 280
rect -45 246 -29 280
rect -129 230 -29 246
rect 29 280 129 318
rect 29 246 45 280
rect 113 246 129 280
rect 29 230 129 246
rect 187 280 287 318
rect 187 246 203 280
rect 271 246 287 280
rect 187 230 287 246
rect 345 280 445 318
rect 345 246 361 280
rect 429 246 445 280
rect 345 230 445 246
rect 503 280 603 318
rect 503 246 519 280
rect 587 246 603 280
rect 503 230 603 246
rect 661 280 761 318
rect 661 246 677 280
rect 745 246 761 280
rect 661 230 761 246
rect 819 280 919 318
rect 819 246 835 280
rect 903 246 919 280
rect 819 230 919 246
rect 977 280 1077 318
rect 977 246 993 280
rect 1061 246 1077 280
rect 977 230 1077 246
rect 1135 280 1235 318
rect 1135 246 1151 280
rect 1219 246 1235 280
rect 1135 230 1235 246
rect 1293 280 1393 318
rect 1293 246 1309 280
rect 1377 246 1393 280
rect 1293 230 1393 246
rect 1451 280 1551 318
rect 1451 246 1467 280
rect 1535 246 1551 280
rect 1451 230 1551 246
rect 1609 280 1709 318
rect 1609 246 1625 280
rect 1693 246 1709 280
rect 1609 230 1709 246
rect 1767 280 1867 318
rect 1767 246 1783 280
rect 1851 246 1867 280
rect 1767 230 1867 246
rect 1925 280 2025 318
rect 1925 246 1941 280
rect 2009 246 2025 280
rect 1925 230 2025 246
rect 2083 280 2183 318
rect 2083 246 2099 280
rect 2167 246 2183 280
rect 2083 230 2183 246
rect 2241 280 2341 318
rect 2241 246 2257 280
rect 2325 246 2341 280
rect 2241 230 2341 246
rect 2399 280 2499 318
rect 2399 246 2415 280
rect 2483 246 2499 280
rect 2399 230 2499 246
rect 2557 280 2657 318
rect 2557 246 2573 280
rect 2641 246 2657 280
rect 2557 230 2657 246
rect 2715 280 2815 318
rect 2715 246 2731 280
rect 2799 246 2815 280
rect 2715 230 2815 246
rect 2873 280 2973 318
rect 2873 246 2889 280
rect 2957 246 2973 280
rect 2873 230 2973 246
rect 3031 280 3131 318
rect 3031 246 3047 280
rect 3115 246 3131 280
rect 3031 230 3131 246
rect -3131 172 -3031 188
rect -3131 138 -3115 172
rect -3047 138 -3031 172
rect -3131 100 -3031 138
rect -2973 172 -2873 188
rect -2973 138 -2957 172
rect -2889 138 -2873 172
rect -2973 100 -2873 138
rect -2815 172 -2715 188
rect -2815 138 -2799 172
rect -2731 138 -2715 172
rect -2815 100 -2715 138
rect -2657 172 -2557 188
rect -2657 138 -2641 172
rect -2573 138 -2557 172
rect -2657 100 -2557 138
rect -2499 172 -2399 188
rect -2499 138 -2483 172
rect -2415 138 -2399 172
rect -2499 100 -2399 138
rect -2341 172 -2241 188
rect -2341 138 -2325 172
rect -2257 138 -2241 172
rect -2341 100 -2241 138
rect -2183 172 -2083 188
rect -2183 138 -2167 172
rect -2099 138 -2083 172
rect -2183 100 -2083 138
rect -2025 172 -1925 188
rect -2025 138 -2009 172
rect -1941 138 -1925 172
rect -2025 100 -1925 138
rect -1867 172 -1767 188
rect -1867 138 -1851 172
rect -1783 138 -1767 172
rect -1867 100 -1767 138
rect -1709 172 -1609 188
rect -1709 138 -1693 172
rect -1625 138 -1609 172
rect -1709 100 -1609 138
rect -1551 172 -1451 188
rect -1551 138 -1535 172
rect -1467 138 -1451 172
rect -1551 100 -1451 138
rect -1393 172 -1293 188
rect -1393 138 -1377 172
rect -1309 138 -1293 172
rect -1393 100 -1293 138
rect -1235 172 -1135 188
rect -1235 138 -1219 172
rect -1151 138 -1135 172
rect -1235 100 -1135 138
rect -1077 172 -977 188
rect -1077 138 -1061 172
rect -993 138 -977 172
rect -1077 100 -977 138
rect -919 172 -819 188
rect -919 138 -903 172
rect -835 138 -819 172
rect -919 100 -819 138
rect -761 172 -661 188
rect -761 138 -745 172
rect -677 138 -661 172
rect -761 100 -661 138
rect -603 172 -503 188
rect -603 138 -587 172
rect -519 138 -503 172
rect -603 100 -503 138
rect -445 172 -345 188
rect -445 138 -429 172
rect -361 138 -345 172
rect -445 100 -345 138
rect -287 172 -187 188
rect -287 138 -271 172
rect -203 138 -187 172
rect -287 100 -187 138
rect -129 172 -29 188
rect -129 138 -113 172
rect -45 138 -29 172
rect -129 100 -29 138
rect 29 172 129 188
rect 29 138 45 172
rect 113 138 129 172
rect 29 100 129 138
rect 187 172 287 188
rect 187 138 203 172
rect 271 138 287 172
rect 187 100 287 138
rect 345 172 445 188
rect 345 138 361 172
rect 429 138 445 172
rect 345 100 445 138
rect 503 172 603 188
rect 503 138 519 172
rect 587 138 603 172
rect 503 100 603 138
rect 661 172 761 188
rect 661 138 677 172
rect 745 138 761 172
rect 661 100 761 138
rect 819 172 919 188
rect 819 138 835 172
rect 903 138 919 172
rect 819 100 919 138
rect 977 172 1077 188
rect 977 138 993 172
rect 1061 138 1077 172
rect 977 100 1077 138
rect 1135 172 1235 188
rect 1135 138 1151 172
rect 1219 138 1235 172
rect 1135 100 1235 138
rect 1293 172 1393 188
rect 1293 138 1309 172
rect 1377 138 1393 172
rect 1293 100 1393 138
rect 1451 172 1551 188
rect 1451 138 1467 172
rect 1535 138 1551 172
rect 1451 100 1551 138
rect 1609 172 1709 188
rect 1609 138 1625 172
rect 1693 138 1709 172
rect 1609 100 1709 138
rect 1767 172 1867 188
rect 1767 138 1783 172
rect 1851 138 1867 172
rect 1767 100 1867 138
rect 1925 172 2025 188
rect 1925 138 1941 172
rect 2009 138 2025 172
rect 1925 100 2025 138
rect 2083 172 2183 188
rect 2083 138 2099 172
rect 2167 138 2183 172
rect 2083 100 2183 138
rect 2241 172 2341 188
rect 2241 138 2257 172
rect 2325 138 2341 172
rect 2241 100 2341 138
rect 2399 172 2499 188
rect 2399 138 2415 172
rect 2483 138 2499 172
rect 2399 100 2499 138
rect 2557 172 2657 188
rect 2557 138 2573 172
rect 2641 138 2657 172
rect 2557 100 2657 138
rect 2715 172 2815 188
rect 2715 138 2731 172
rect 2799 138 2815 172
rect 2715 100 2815 138
rect 2873 172 2973 188
rect 2873 138 2889 172
rect 2957 138 2973 172
rect 2873 100 2973 138
rect 3031 172 3131 188
rect 3031 138 3047 172
rect 3115 138 3131 172
rect 3031 100 3131 138
rect -3131 -138 -3031 -100
rect -3131 -172 -3115 -138
rect -3047 -172 -3031 -138
rect -3131 -188 -3031 -172
rect -2973 -138 -2873 -100
rect -2973 -172 -2957 -138
rect -2889 -172 -2873 -138
rect -2973 -188 -2873 -172
rect -2815 -138 -2715 -100
rect -2815 -172 -2799 -138
rect -2731 -172 -2715 -138
rect -2815 -188 -2715 -172
rect -2657 -138 -2557 -100
rect -2657 -172 -2641 -138
rect -2573 -172 -2557 -138
rect -2657 -188 -2557 -172
rect -2499 -138 -2399 -100
rect -2499 -172 -2483 -138
rect -2415 -172 -2399 -138
rect -2499 -188 -2399 -172
rect -2341 -138 -2241 -100
rect -2341 -172 -2325 -138
rect -2257 -172 -2241 -138
rect -2341 -188 -2241 -172
rect -2183 -138 -2083 -100
rect -2183 -172 -2167 -138
rect -2099 -172 -2083 -138
rect -2183 -188 -2083 -172
rect -2025 -138 -1925 -100
rect -2025 -172 -2009 -138
rect -1941 -172 -1925 -138
rect -2025 -188 -1925 -172
rect -1867 -138 -1767 -100
rect -1867 -172 -1851 -138
rect -1783 -172 -1767 -138
rect -1867 -188 -1767 -172
rect -1709 -138 -1609 -100
rect -1709 -172 -1693 -138
rect -1625 -172 -1609 -138
rect -1709 -188 -1609 -172
rect -1551 -138 -1451 -100
rect -1551 -172 -1535 -138
rect -1467 -172 -1451 -138
rect -1551 -188 -1451 -172
rect -1393 -138 -1293 -100
rect -1393 -172 -1377 -138
rect -1309 -172 -1293 -138
rect -1393 -188 -1293 -172
rect -1235 -138 -1135 -100
rect -1235 -172 -1219 -138
rect -1151 -172 -1135 -138
rect -1235 -188 -1135 -172
rect -1077 -138 -977 -100
rect -1077 -172 -1061 -138
rect -993 -172 -977 -138
rect -1077 -188 -977 -172
rect -919 -138 -819 -100
rect -919 -172 -903 -138
rect -835 -172 -819 -138
rect -919 -188 -819 -172
rect -761 -138 -661 -100
rect -761 -172 -745 -138
rect -677 -172 -661 -138
rect -761 -188 -661 -172
rect -603 -138 -503 -100
rect -603 -172 -587 -138
rect -519 -172 -503 -138
rect -603 -188 -503 -172
rect -445 -138 -345 -100
rect -445 -172 -429 -138
rect -361 -172 -345 -138
rect -445 -188 -345 -172
rect -287 -138 -187 -100
rect -287 -172 -271 -138
rect -203 -172 -187 -138
rect -287 -188 -187 -172
rect -129 -138 -29 -100
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect -129 -188 -29 -172
rect 29 -138 129 -100
rect 29 -172 45 -138
rect 113 -172 129 -138
rect 29 -188 129 -172
rect 187 -138 287 -100
rect 187 -172 203 -138
rect 271 -172 287 -138
rect 187 -188 287 -172
rect 345 -138 445 -100
rect 345 -172 361 -138
rect 429 -172 445 -138
rect 345 -188 445 -172
rect 503 -138 603 -100
rect 503 -172 519 -138
rect 587 -172 603 -138
rect 503 -188 603 -172
rect 661 -138 761 -100
rect 661 -172 677 -138
rect 745 -172 761 -138
rect 661 -188 761 -172
rect 819 -138 919 -100
rect 819 -172 835 -138
rect 903 -172 919 -138
rect 819 -188 919 -172
rect 977 -138 1077 -100
rect 977 -172 993 -138
rect 1061 -172 1077 -138
rect 977 -188 1077 -172
rect 1135 -138 1235 -100
rect 1135 -172 1151 -138
rect 1219 -172 1235 -138
rect 1135 -188 1235 -172
rect 1293 -138 1393 -100
rect 1293 -172 1309 -138
rect 1377 -172 1393 -138
rect 1293 -188 1393 -172
rect 1451 -138 1551 -100
rect 1451 -172 1467 -138
rect 1535 -172 1551 -138
rect 1451 -188 1551 -172
rect 1609 -138 1709 -100
rect 1609 -172 1625 -138
rect 1693 -172 1709 -138
rect 1609 -188 1709 -172
rect 1767 -138 1867 -100
rect 1767 -172 1783 -138
rect 1851 -172 1867 -138
rect 1767 -188 1867 -172
rect 1925 -138 2025 -100
rect 1925 -172 1941 -138
rect 2009 -172 2025 -138
rect 1925 -188 2025 -172
rect 2083 -138 2183 -100
rect 2083 -172 2099 -138
rect 2167 -172 2183 -138
rect 2083 -188 2183 -172
rect 2241 -138 2341 -100
rect 2241 -172 2257 -138
rect 2325 -172 2341 -138
rect 2241 -188 2341 -172
rect 2399 -138 2499 -100
rect 2399 -172 2415 -138
rect 2483 -172 2499 -138
rect 2399 -188 2499 -172
rect 2557 -138 2657 -100
rect 2557 -172 2573 -138
rect 2641 -172 2657 -138
rect 2557 -188 2657 -172
rect 2715 -138 2815 -100
rect 2715 -172 2731 -138
rect 2799 -172 2815 -138
rect 2715 -188 2815 -172
rect 2873 -138 2973 -100
rect 2873 -172 2889 -138
rect 2957 -172 2973 -138
rect 2873 -188 2973 -172
rect 3031 -138 3131 -100
rect 3031 -172 3047 -138
rect 3115 -172 3131 -138
rect 3031 -188 3131 -172
rect -3131 -246 -3031 -230
rect -3131 -280 -3115 -246
rect -3047 -280 -3031 -246
rect -3131 -318 -3031 -280
rect -2973 -246 -2873 -230
rect -2973 -280 -2957 -246
rect -2889 -280 -2873 -246
rect -2973 -318 -2873 -280
rect -2815 -246 -2715 -230
rect -2815 -280 -2799 -246
rect -2731 -280 -2715 -246
rect -2815 -318 -2715 -280
rect -2657 -246 -2557 -230
rect -2657 -280 -2641 -246
rect -2573 -280 -2557 -246
rect -2657 -318 -2557 -280
rect -2499 -246 -2399 -230
rect -2499 -280 -2483 -246
rect -2415 -280 -2399 -246
rect -2499 -318 -2399 -280
rect -2341 -246 -2241 -230
rect -2341 -280 -2325 -246
rect -2257 -280 -2241 -246
rect -2341 -318 -2241 -280
rect -2183 -246 -2083 -230
rect -2183 -280 -2167 -246
rect -2099 -280 -2083 -246
rect -2183 -318 -2083 -280
rect -2025 -246 -1925 -230
rect -2025 -280 -2009 -246
rect -1941 -280 -1925 -246
rect -2025 -318 -1925 -280
rect -1867 -246 -1767 -230
rect -1867 -280 -1851 -246
rect -1783 -280 -1767 -246
rect -1867 -318 -1767 -280
rect -1709 -246 -1609 -230
rect -1709 -280 -1693 -246
rect -1625 -280 -1609 -246
rect -1709 -318 -1609 -280
rect -1551 -246 -1451 -230
rect -1551 -280 -1535 -246
rect -1467 -280 -1451 -246
rect -1551 -318 -1451 -280
rect -1393 -246 -1293 -230
rect -1393 -280 -1377 -246
rect -1309 -280 -1293 -246
rect -1393 -318 -1293 -280
rect -1235 -246 -1135 -230
rect -1235 -280 -1219 -246
rect -1151 -280 -1135 -246
rect -1235 -318 -1135 -280
rect -1077 -246 -977 -230
rect -1077 -280 -1061 -246
rect -993 -280 -977 -246
rect -1077 -318 -977 -280
rect -919 -246 -819 -230
rect -919 -280 -903 -246
rect -835 -280 -819 -246
rect -919 -318 -819 -280
rect -761 -246 -661 -230
rect -761 -280 -745 -246
rect -677 -280 -661 -246
rect -761 -318 -661 -280
rect -603 -246 -503 -230
rect -603 -280 -587 -246
rect -519 -280 -503 -246
rect -603 -318 -503 -280
rect -445 -246 -345 -230
rect -445 -280 -429 -246
rect -361 -280 -345 -246
rect -445 -318 -345 -280
rect -287 -246 -187 -230
rect -287 -280 -271 -246
rect -203 -280 -187 -246
rect -287 -318 -187 -280
rect -129 -246 -29 -230
rect -129 -280 -113 -246
rect -45 -280 -29 -246
rect -129 -318 -29 -280
rect 29 -246 129 -230
rect 29 -280 45 -246
rect 113 -280 129 -246
rect 29 -318 129 -280
rect 187 -246 287 -230
rect 187 -280 203 -246
rect 271 -280 287 -246
rect 187 -318 287 -280
rect 345 -246 445 -230
rect 345 -280 361 -246
rect 429 -280 445 -246
rect 345 -318 445 -280
rect 503 -246 603 -230
rect 503 -280 519 -246
rect 587 -280 603 -246
rect 503 -318 603 -280
rect 661 -246 761 -230
rect 661 -280 677 -246
rect 745 -280 761 -246
rect 661 -318 761 -280
rect 819 -246 919 -230
rect 819 -280 835 -246
rect 903 -280 919 -246
rect 819 -318 919 -280
rect 977 -246 1077 -230
rect 977 -280 993 -246
rect 1061 -280 1077 -246
rect 977 -318 1077 -280
rect 1135 -246 1235 -230
rect 1135 -280 1151 -246
rect 1219 -280 1235 -246
rect 1135 -318 1235 -280
rect 1293 -246 1393 -230
rect 1293 -280 1309 -246
rect 1377 -280 1393 -246
rect 1293 -318 1393 -280
rect 1451 -246 1551 -230
rect 1451 -280 1467 -246
rect 1535 -280 1551 -246
rect 1451 -318 1551 -280
rect 1609 -246 1709 -230
rect 1609 -280 1625 -246
rect 1693 -280 1709 -246
rect 1609 -318 1709 -280
rect 1767 -246 1867 -230
rect 1767 -280 1783 -246
rect 1851 -280 1867 -246
rect 1767 -318 1867 -280
rect 1925 -246 2025 -230
rect 1925 -280 1941 -246
rect 2009 -280 2025 -246
rect 1925 -318 2025 -280
rect 2083 -246 2183 -230
rect 2083 -280 2099 -246
rect 2167 -280 2183 -246
rect 2083 -318 2183 -280
rect 2241 -246 2341 -230
rect 2241 -280 2257 -246
rect 2325 -280 2341 -246
rect 2241 -318 2341 -280
rect 2399 -246 2499 -230
rect 2399 -280 2415 -246
rect 2483 -280 2499 -246
rect 2399 -318 2499 -280
rect 2557 -246 2657 -230
rect 2557 -280 2573 -246
rect 2641 -280 2657 -246
rect 2557 -318 2657 -280
rect 2715 -246 2815 -230
rect 2715 -280 2731 -246
rect 2799 -280 2815 -246
rect 2715 -318 2815 -280
rect 2873 -246 2973 -230
rect 2873 -280 2889 -246
rect 2957 -280 2973 -246
rect 2873 -318 2973 -280
rect 3031 -246 3131 -230
rect 3031 -280 3047 -246
rect 3115 -280 3131 -246
rect 3031 -318 3131 -280
rect -3131 -556 -3031 -518
rect -3131 -590 -3115 -556
rect -3047 -590 -3031 -556
rect -3131 -606 -3031 -590
rect -2973 -556 -2873 -518
rect -2973 -590 -2957 -556
rect -2889 -590 -2873 -556
rect -2973 -606 -2873 -590
rect -2815 -556 -2715 -518
rect -2815 -590 -2799 -556
rect -2731 -590 -2715 -556
rect -2815 -606 -2715 -590
rect -2657 -556 -2557 -518
rect -2657 -590 -2641 -556
rect -2573 -590 -2557 -556
rect -2657 -606 -2557 -590
rect -2499 -556 -2399 -518
rect -2499 -590 -2483 -556
rect -2415 -590 -2399 -556
rect -2499 -606 -2399 -590
rect -2341 -556 -2241 -518
rect -2341 -590 -2325 -556
rect -2257 -590 -2241 -556
rect -2341 -606 -2241 -590
rect -2183 -556 -2083 -518
rect -2183 -590 -2167 -556
rect -2099 -590 -2083 -556
rect -2183 -606 -2083 -590
rect -2025 -556 -1925 -518
rect -2025 -590 -2009 -556
rect -1941 -590 -1925 -556
rect -2025 -606 -1925 -590
rect -1867 -556 -1767 -518
rect -1867 -590 -1851 -556
rect -1783 -590 -1767 -556
rect -1867 -606 -1767 -590
rect -1709 -556 -1609 -518
rect -1709 -590 -1693 -556
rect -1625 -590 -1609 -556
rect -1709 -606 -1609 -590
rect -1551 -556 -1451 -518
rect -1551 -590 -1535 -556
rect -1467 -590 -1451 -556
rect -1551 -606 -1451 -590
rect -1393 -556 -1293 -518
rect -1393 -590 -1377 -556
rect -1309 -590 -1293 -556
rect -1393 -606 -1293 -590
rect -1235 -556 -1135 -518
rect -1235 -590 -1219 -556
rect -1151 -590 -1135 -556
rect -1235 -606 -1135 -590
rect -1077 -556 -977 -518
rect -1077 -590 -1061 -556
rect -993 -590 -977 -556
rect -1077 -606 -977 -590
rect -919 -556 -819 -518
rect -919 -590 -903 -556
rect -835 -590 -819 -556
rect -919 -606 -819 -590
rect -761 -556 -661 -518
rect -761 -590 -745 -556
rect -677 -590 -661 -556
rect -761 -606 -661 -590
rect -603 -556 -503 -518
rect -603 -590 -587 -556
rect -519 -590 -503 -556
rect -603 -606 -503 -590
rect -445 -556 -345 -518
rect -445 -590 -429 -556
rect -361 -590 -345 -556
rect -445 -606 -345 -590
rect -287 -556 -187 -518
rect -287 -590 -271 -556
rect -203 -590 -187 -556
rect -287 -606 -187 -590
rect -129 -556 -29 -518
rect -129 -590 -113 -556
rect -45 -590 -29 -556
rect -129 -606 -29 -590
rect 29 -556 129 -518
rect 29 -590 45 -556
rect 113 -590 129 -556
rect 29 -606 129 -590
rect 187 -556 287 -518
rect 187 -590 203 -556
rect 271 -590 287 -556
rect 187 -606 287 -590
rect 345 -556 445 -518
rect 345 -590 361 -556
rect 429 -590 445 -556
rect 345 -606 445 -590
rect 503 -556 603 -518
rect 503 -590 519 -556
rect 587 -590 603 -556
rect 503 -606 603 -590
rect 661 -556 761 -518
rect 661 -590 677 -556
rect 745 -590 761 -556
rect 661 -606 761 -590
rect 819 -556 919 -518
rect 819 -590 835 -556
rect 903 -590 919 -556
rect 819 -606 919 -590
rect 977 -556 1077 -518
rect 977 -590 993 -556
rect 1061 -590 1077 -556
rect 977 -606 1077 -590
rect 1135 -556 1235 -518
rect 1135 -590 1151 -556
rect 1219 -590 1235 -556
rect 1135 -606 1235 -590
rect 1293 -556 1393 -518
rect 1293 -590 1309 -556
rect 1377 -590 1393 -556
rect 1293 -606 1393 -590
rect 1451 -556 1551 -518
rect 1451 -590 1467 -556
rect 1535 -590 1551 -556
rect 1451 -606 1551 -590
rect 1609 -556 1709 -518
rect 1609 -590 1625 -556
rect 1693 -590 1709 -556
rect 1609 -606 1709 -590
rect 1767 -556 1867 -518
rect 1767 -590 1783 -556
rect 1851 -590 1867 -556
rect 1767 -606 1867 -590
rect 1925 -556 2025 -518
rect 1925 -590 1941 -556
rect 2009 -590 2025 -556
rect 1925 -606 2025 -590
rect 2083 -556 2183 -518
rect 2083 -590 2099 -556
rect 2167 -590 2183 -556
rect 2083 -606 2183 -590
rect 2241 -556 2341 -518
rect 2241 -590 2257 -556
rect 2325 -590 2341 -556
rect 2241 -606 2341 -590
rect 2399 -556 2499 -518
rect 2399 -590 2415 -556
rect 2483 -590 2499 -556
rect 2399 -606 2499 -590
rect 2557 -556 2657 -518
rect 2557 -590 2573 -556
rect 2641 -590 2657 -556
rect 2557 -606 2657 -590
rect 2715 -556 2815 -518
rect 2715 -590 2731 -556
rect 2799 -590 2815 -556
rect 2715 -606 2815 -590
rect 2873 -556 2973 -518
rect 2873 -590 2889 -556
rect 2957 -590 2973 -556
rect 2873 -606 2973 -590
rect 3031 -556 3131 -518
rect 3031 -590 3047 -556
rect 3115 -590 3131 -556
rect 3031 -606 3131 -590
<< polycont >>
rect -3115 556 -3047 590
rect -2957 556 -2889 590
rect -2799 556 -2731 590
rect -2641 556 -2573 590
rect -2483 556 -2415 590
rect -2325 556 -2257 590
rect -2167 556 -2099 590
rect -2009 556 -1941 590
rect -1851 556 -1783 590
rect -1693 556 -1625 590
rect -1535 556 -1467 590
rect -1377 556 -1309 590
rect -1219 556 -1151 590
rect -1061 556 -993 590
rect -903 556 -835 590
rect -745 556 -677 590
rect -587 556 -519 590
rect -429 556 -361 590
rect -271 556 -203 590
rect -113 556 -45 590
rect 45 556 113 590
rect 203 556 271 590
rect 361 556 429 590
rect 519 556 587 590
rect 677 556 745 590
rect 835 556 903 590
rect 993 556 1061 590
rect 1151 556 1219 590
rect 1309 556 1377 590
rect 1467 556 1535 590
rect 1625 556 1693 590
rect 1783 556 1851 590
rect 1941 556 2009 590
rect 2099 556 2167 590
rect 2257 556 2325 590
rect 2415 556 2483 590
rect 2573 556 2641 590
rect 2731 556 2799 590
rect 2889 556 2957 590
rect 3047 556 3115 590
rect -3115 246 -3047 280
rect -2957 246 -2889 280
rect -2799 246 -2731 280
rect -2641 246 -2573 280
rect -2483 246 -2415 280
rect -2325 246 -2257 280
rect -2167 246 -2099 280
rect -2009 246 -1941 280
rect -1851 246 -1783 280
rect -1693 246 -1625 280
rect -1535 246 -1467 280
rect -1377 246 -1309 280
rect -1219 246 -1151 280
rect -1061 246 -993 280
rect -903 246 -835 280
rect -745 246 -677 280
rect -587 246 -519 280
rect -429 246 -361 280
rect -271 246 -203 280
rect -113 246 -45 280
rect 45 246 113 280
rect 203 246 271 280
rect 361 246 429 280
rect 519 246 587 280
rect 677 246 745 280
rect 835 246 903 280
rect 993 246 1061 280
rect 1151 246 1219 280
rect 1309 246 1377 280
rect 1467 246 1535 280
rect 1625 246 1693 280
rect 1783 246 1851 280
rect 1941 246 2009 280
rect 2099 246 2167 280
rect 2257 246 2325 280
rect 2415 246 2483 280
rect 2573 246 2641 280
rect 2731 246 2799 280
rect 2889 246 2957 280
rect 3047 246 3115 280
rect -3115 138 -3047 172
rect -2957 138 -2889 172
rect -2799 138 -2731 172
rect -2641 138 -2573 172
rect -2483 138 -2415 172
rect -2325 138 -2257 172
rect -2167 138 -2099 172
rect -2009 138 -1941 172
rect -1851 138 -1783 172
rect -1693 138 -1625 172
rect -1535 138 -1467 172
rect -1377 138 -1309 172
rect -1219 138 -1151 172
rect -1061 138 -993 172
rect -903 138 -835 172
rect -745 138 -677 172
rect -587 138 -519 172
rect -429 138 -361 172
rect -271 138 -203 172
rect -113 138 -45 172
rect 45 138 113 172
rect 203 138 271 172
rect 361 138 429 172
rect 519 138 587 172
rect 677 138 745 172
rect 835 138 903 172
rect 993 138 1061 172
rect 1151 138 1219 172
rect 1309 138 1377 172
rect 1467 138 1535 172
rect 1625 138 1693 172
rect 1783 138 1851 172
rect 1941 138 2009 172
rect 2099 138 2167 172
rect 2257 138 2325 172
rect 2415 138 2483 172
rect 2573 138 2641 172
rect 2731 138 2799 172
rect 2889 138 2957 172
rect 3047 138 3115 172
rect -3115 -172 -3047 -138
rect -2957 -172 -2889 -138
rect -2799 -172 -2731 -138
rect -2641 -172 -2573 -138
rect -2483 -172 -2415 -138
rect -2325 -172 -2257 -138
rect -2167 -172 -2099 -138
rect -2009 -172 -1941 -138
rect -1851 -172 -1783 -138
rect -1693 -172 -1625 -138
rect -1535 -172 -1467 -138
rect -1377 -172 -1309 -138
rect -1219 -172 -1151 -138
rect -1061 -172 -993 -138
rect -903 -172 -835 -138
rect -745 -172 -677 -138
rect -587 -172 -519 -138
rect -429 -172 -361 -138
rect -271 -172 -203 -138
rect -113 -172 -45 -138
rect 45 -172 113 -138
rect 203 -172 271 -138
rect 361 -172 429 -138
rect 519 -172 587 -138
rect 677 -172 745 -138
rect 835 -172 903 -138
rect 993 -172 1061 -138
rect 1151 -172 1219 -138
rect 1309 -172 1377 -138
rect 1467 -172 1535 -138
rect 1625 -172 1693 -138
rect 1783 -172 1851 -138
rect 1941 -172 2009 -138
rect 2099 -172 2167 -138
rect 2257 -172 2325 -138
rect 2415 -172 2483 -138
rect 2573 -172 2641 -138
rect 2731 -172 2799 -138
rect 2889 -172 2957 -138
rect 3047 -172 3115 -138
rect -3115 -280 -3047 -246
rect -2957 -280 -2889 -246
rect -2799 -280 -2731 -246
rect -2641 -280 -2573 -246
rect -2483 -280 -2415 -246
rect -2325 -280 -2257 -246
rect -2167 -280 -2099 -246
rect -2009 -280 -1941 -246
rect -1851 -280 -1783 -246
rect -1693 -280 -1625 -246
rect -1535 -280 -1467 -246
rect -1377 -280 -1309 -246
rect -1219 -280 -1151 -246
rect -1061 -280 -993 -246
rect -903 -280 -835 -246
rect -745 -280 -677 -246
rect -587 -280 -519 -246
rect -429 -280 -361 -246
rect -271 -280 -203 -246
rect -113 -280 -45 -246
rect 45 -280 113 -246
rect 203 -280 271 -246
rect 361 -280 429 -246
rect 519 -280 587 -246
rect 677 -280 745 -246
rect 835 -280 903 -246
rect 993 -280 1061 -246
rect 1151 -280 1219 -246
rect 1309 -280 1377 -246
rect 1467 -280 1535 -246
rect 1625 -280 1693 -246
rect 1783 -280 1851 -246
rect 1941 -280 2009 -246
rect 2099 -280 2167 -246
rect 2257 -280 2325 -246
rect 2415 -280 2483 -246
rect 2573 -280 2641 -246
rect 2731 -280 2799 -246
rect 2889 -280 2957 -246
rect 3047 -280 3115 -246
rect -3115 -590 -3047 -556
rect -2957 -590 -2889 -556
rect -2799 -590 -2731 -556
rect -2641 -590 -2573 -556
rect -2483 -590 -2415 -556
rect -2325 -590 -2257 -556
rect -2167 -590 -2099 -556
rect -2009 -590 -1941 -556
rect -1851 -590 -1783 -556
rect -1693 -590 -1625 -556
rect -1535 -590 -1467 -556
rect -1377 -590 -1309 -556
rect -1219 -590 -1151 -556
rect -1061 -590 -993 -556
rect -903 -590 -835 -556
rect -745 -590 -677 -556
rect -587 -590 -519 -556
rect -429 -590 -361 -556
rect -271 -590 -203 -556
rect -113 -590 -45 -556
rect 45 -590 113 -556
rect 203 -590 271 -556
rect 361 -590 429 -556
rect 519 -590 587 -556
rect 677 -590 745 -556
rect 835 -590 903 -556
rect 993 -590 1061 -556
rect 1151 -590 1219 -556
rect 1309 -590 1377 -556
rect 1467 -590 1535 -556
rect 1625 -590 1693 -556
rect 1783 -590 1851 -556
rect 1941 -590 2009 -556
rect 2099 -590 2167 -556
rect 2257 -590 2325 -556
rect 2415 -590 2483 -556
rect 2573 -590 2641 -556
rect 2731 -590 2799 -556
rect 2889 -590 2957 -556
rect 3047 -590 3115 -556
<< locali >>
rect -3311 694 -3215 728
rect 3215 694 3311 728
rect -3311 632 -3277 694
rect 3277 632 3311 694
rect -3131 556 -3115 590
rect -3047 556 -3031 590
rect -2973 556 -2957 590
rect -2889 556 -2873 590
rect -2815 556 -2799 590
rect -2731 556 -2715 590
rect -2657 556 -2641 590
rect -2573 556 -2557 590
rect -2499 556 -2483 590
rect -2415 556 -2399 590
rect -2341 556 -2325 590
rect -2257 556 -2241 590
rect -2183 556 -2167 590
rect -2099 556 -2083 590
rect -2025 556 -2009 590
rect -1941 556 -1925 590
rect -1867 556 -1851 590
rect -1783 556 -1767 590
rect -1709 556 -1693 590
rect -1625 556 -1609 590
rect -1551 556 -1535 590
rect -1467 556 -1451 590
rect -1393 556 -1377 590
rect -1309 556 -1293 590
rect -1235 556 -1219 590
rect -1151 556 -1135 590
rect -1077 556 -1061 590
rect -993 556 -977 590
rect -919 556 -903 590
rect -835 556 -819 590
rect -761 556 -745 590
rect -677 556 -661 590
rect -603 556 -587 590
rect -519 556 -503 590
rect -445 556 -429 590
rect -361 556 -345 590
rect -287 556 -271 590
rect -203 556 -187 590
rect -129 556 -113 590
rect -45 556 -29 590
rect 29 556 45 590
rect 113 556 129 590
rect 187 556 203 590
rect 271 556 287 590
rect 345 556 361 590
rect 429 556 445 590
rect 503 556 519 590
rect 587 556 603 590
rect 661 556 677 590
rect 745 556 761 590
rect 819 556 835 590
rect 903 556 919 590
rect 977 556 993 590
rect 1061 556 1077 590
rect 1135 556 1151 590
rect 1219 556 1235 590
rect 1293 556 1309 590
rect 1377 556 1393 590
rect 1451 556 1467 590
rect 1535 556 1551 590
rect 1609 556 1625 590
rect 1693 556 1709 590
rect 1767 556 1783 590
rect 1851 556 1867 590
rect 1925 556 1941 590
rect 2009 556 2025 590
rect 2083 556 2099 590
rect 2167 556 2183 590
rect 2241 556 2257 590
rect 2325 556 2341 590
rect 2399 556 2415 590
rect 2483 556 2499 590
rect 2557 556 2573 590
rect 2641 556 2657 590
rect 2715 556 2731 590
rect 2799 556 2815 590
rect 2873 556 2889 590
rect 2957 556 2973 590
rect 3031 556 3047 590
rect 3115 556 3131 590
rect -3177 506 -3143 522
rect -3177 314 -3143 330
rect -3019 506 -2985 522
rect -3019 314 -2985 330
rect -2861 506 -2827 522
rect -2861 314 -2827 330
rect -2703 506 -2669 522
rect -2703 314 -2669 330
rect -2545 506 -2511 522
rect -2545 314 -2511 330
rect -2387 506 -2353 522
rect -2387 314 -2353 330
rect -2229 506 -2195 522
rect -2229 314 -2195 330
rect -2071 506 -2037 522
rect -2071 314 -2037 330
rect -1913 506 -1879 522
rect -1913 314 -1879 330
rect -1755 506 -1721 522
rect -1755 314 -1721 330
rect -1597 506 -1563 522
rect -1597 314 -1563 330
rect -1439 506 -1405 522
rect -1439 314 -1405 330
rect -1281 506 -1247 522
rect -1281 314 -1247 330
rect -1123 506 -1089 522
rect -1123 314 -1089 330
rect -965 506 -931 522
rect -965 314 -931 330
rect -807 506 -773 522
rect -807 314 -773 330
rect -649 506 -615 522
rect -649 314 -615 330
rect -491 506 -457 522
rect -491 314 -457 330
rect -333 506 -299 522
rect -333 314 -299 330
rect -175 506 -141 522
rect -175 314 -141 330
rect -17 506 17 522
rect -17 314 17 330
rect 141 506 175 522
rect 141 314 175 330
rect 299 506 333 522
rect 299 314 333 330
rect 457 506 491 522
rect 457 314 491 330
rect 615 506 649 522
rect 615 314 649 330
rect 773 506 807 522
rect 773 314 807 330
rect 931 506 965 522
rect 931 314 965 330
rect 1089 506 1123 522
rect 1089 314 1123 330
rect 1247 506 1281 522
rect 1247 314 1281 330
rect 1405 506 1439 522
rect 1405 314 1439 330
rect 1563 506 1597 522
rect 1563 314 1597 330
rect 1721 506 1755 522
rect 1721 314 1755 330
rect 1879 506 1913 522
rect 1879 314 1913 330
rect 2037 506 2071 522
rect 2037 314 2071 330
rect 2195 506 2229 522
rect 2195 314 2229 330
rect 2353 506 2387 522
rect 2353 314 2387 330
rect 2511 506 2545 522
rect 2511 314 2545 330
rect 2669 506 2703 522
rect 2669 314 2703 330
rect 2827 506 2861 522
rect 2827 314 2861 330
rect 2985 506 3019 522
rect 2985 314 3019 330
rect 3143 506 3177 522
rect 3143 314 3177 330
rect -3131 246 -3115 280
rect -3047 246 -3031 280
rect -2973 246 -2957 280
rect -2889 246 -2873 280
rect -2815 246 -2799 280
rect -2731 246 -2715 280
rect -2657 246 -2641 280
rect -2573 246 -2557 280
rect -2499 246 -2483 280
rect -2415 246 -2399 280
rect -2341 246 -2325 280
rect -2257 246 -2241 280
rect -2183 246 -2167 280
rect -2099 246 -2083 280
rect -2025 246 -2009 280
rect -1941 246 -1925 280
rect -1867 246 -1851 280
rect -1783 246 -1767 280
rect -1709 246 -1693 280
rect -1625 246 -1609 280
rect -1551 246 -1535 280
rect -1467 246 -1451 280
rect -1393 246 -1377 280
rect -1309 246 -1293 280
rect -1235 246 -1219 280
rect -1151 246 -1135 280
rect -1077 246 -1061 280
rect -993 246 -977 280
rect -919 246 -903 280
rect -835 246 -819 280
rect -761 246 -745 280
rect -677 246 -661 280
rect -603 246 -587 280
rect -519 246 -503 280
rect -445 246 -429 280
rect -361 246 -345 280
rect -287 246 -271 280
rect -203 246 -187 280
rect -129 246 -113 280
rect -45 246 -29 280
rect 29 246 45 280
rect 113 246 129 280
rect 187 246 203 280
rect 271 246 287 280
rect 345 246 361 280
rect 429 246 445 280
rect 503 246 519 280
rect 587 246 603 280
rect 661 246 677 280
rect 745 246 761 280
rect 819 246 835 280
rect 903 246 919 280
rect 977 246 993 280
rect 1061 246 1077 280
rect 1135 246 1151 280
rect 1219 246 1235 280
rect 1293 246 1309 280
rect 1377 246 1393 280
rect 1451 246 1467 280
rect 1535 246 1551 280
rect 1609 246 1625 280
rect 1693 246 1709 280
rect 1767 246 1783 280
rect 1851 246 1867 280
rect 1925 246 1941 280
rect 2009 246 2025 280
rect 2083 246 2099 280
rect 2167 246 2183 280
rect 2241 246 2257 280
rect 2325 246 2341 280
rect 2399 246 2415 280
rect 2483 246 2499 280
rect 2557 246 2573 280
rect 2641 246 2657 280
rect 2715 246 2731 280
rect 2799 246 2815 280
rect 2873 246 2889 280
rect 2957 246 2973 280
rect 3031 246 3047 280
rect 3115 246 3131 280
rect -3131 138 -3115 172
rect -3047 138 -3031 172
rect -2973 138 -2957 172
rect -2889 138 -2873 172
rect -2815 138 -2799 172
rect -2731 138 -2715 172
rect -2657 138 -2641 172
rect -2573 138 -2557 172
rect -2499 138 -2483 172
rect -2415 138 -2399 172
rect -2341 138 -2325 172
rect -2257 138 -2241 172
rect -2183 138 -2167 172
rect -2099 138 -2083 172
rect -2025 138 -2009 172
rect -1941 138 -1925 172
rect -1867 138 -1851 172
rect -1783 138 -1767 172
rect -1709 138 -1693 172
rect -1625 138 -1609 172
rect -1551 138 -1535 172
rect -1467 138 -1451 172
rect -1393 138 -1377 172
rect -1309 138 -1293 172
rect -1235 138 -1219 172
rect -1151 138 -1135 172
rect -1077 138 -1061 172
rect -993 138 -977 172
rect -919 138 -903 172
rect -835 138 -819 172
rect -761 138 -745 172
rect -677 138 -661 172
rect -603 138 -587 172
rect -519 138 -503 172
rect -445 138 -429 172
rect -361 138 -345 172
rect -287 138 -271 172
rect -203 138 -187 172
rect -129 138 -113 172
rect -45 138 -29 172
rect 29 138 45 172
rect 113 138 129 172
rect 187 138 203 172
rect 271 138 287 172
rect 345 138 361 172
rect 429 138 445 172
rect 503 138 519 172
rect 587 138 603 172
rect 661 138 677 172
rect 745 138 761 172
rect 819 138 835 172
rect 903 138 919 172
rect 977 138 993 172
rect 1061 138 1077 172
rect 1135 138 1151 172
rect 1219 138 1235 172
rect 1293 138 1309 172
rect 1377 138 1393 172
rect 1451 138 1467 172
rect 1535 138 1551 172
rect 1609 138 1625 172
rect 1693 138 1709 172
rect 1767 138 1783 172
rect 1851 138 1867 172
rect 1925 138 1941 172
rect 2009 138 2025 172
rect 2083 138 2099 172
rect 2167 138 2183 172
rect 2241 138 2257 172
rect 2325 138 2341 172
rect 2399 138 2415 172
rect 2483 138 2499 172
rect 2557 138 2573 172
rect 2641 138 2657 172
rect 2715 138 2731 172
rect 2799 138 2815 172
rect 2873 138 2889 172
rect 2957 138 2973 172
rect 3031 138 3047 172
rect 3115 138 3131 172
rect -3177 88 -3143 104
rect -3177 -104 -3143 -88
rect -3019 88 -2985 104
rect -3019 -104 -2985 -88
rect -2861 88 -2827 104
rect -2861 -104 -2827 -88
rect -2703 88 -2669 104
rect -2703 -104 -2669 -88
rect -2545 88 -2511 104
rect -2545 -104 -2511 -88
rect -2387 88 -2353 104
rect -2387 -104 -2353 -88
rect -2229 88 -2195 104
rect -2229 -104 -2195 -88
rect -2071 88 -2037 104
rect -2071 -104 -2037 -88
rect -1913 88 -1879 104
rect -1913 -104 -1879 -88
rect -1755 88 -1721 104
rect -1755 -104 -1721 -88
rect -1597 88 -1563 104
rect -1597 -104 -1563 -88
rect -1439 88 -1405 104
rect -1439 -104 -1405 -88
rect -1281 88 -1247 104
rect -1281 -104 -1247 -88
rect -1123 88 -1089 104
rect -1123 -104 -1089 -88
rect -965 88 -931 104
rect -965 -104 -931 -88
rect -807 88 -773 104
rect -807 -104 -773 -88
rect -649 88 -615 104
rect -649 -104 -615 -88
rect -491 88 -457 104
rect -491 -104 -457 -88
rect -333 88 -299 104
rect -333 -104 -299 -88
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect 299 88 333 104
rect 299 -104 333 -88
rect 457 88 491 104
rect 457 -104 491 -88
rect 615 88 649 104
rect 615 -104 649 -88
rect 773 88 807 104
rect 773 -104 807 -88
rect 931 88 965 104
rect 931 -104 965 -88
rect 1089 88 1123 104
rect 1089 -104 1123 -88
rect 1247 88 1281 104
rect 1247 -104 1281 -88
rect 1405 88 1439 104
rect 1405 -104 1439 -88
rect 1563 88 1597 104
rect 1563 -104 1597 -88
rect 1721 88 1755 104
rect 1721 -104 1755 -88
rect 1879 88 1913 104
rect 1879 -104 1913 -88
rect 2037 88 2071 104
rect 2037 -104 2071 -88
rect 2195 88 2229 104
rect 2195 -104 2229 -88
rect 2353 88 2387 104
rect 2353 -104 2387 -88
rect 2511 88 2545 104
rect 2511 -104 2545 -88
rect 2669 88 2703 104
rect 2669 -104 2703 -88
rect 2827 88 2861 104
rect 2827 -104 2861 -88
rect 2985 88 3019 104
rect 2985 -104 3019 -88
rect 3143 88 3177 104
rect 3143 -104 3177 -88
rect -3131 -172 -3115 -138
rect -3047 -172 -3031 -138
rect -2973 -172 -2957 -138
rect -2889 -172 -2873 -138
rect -2815 -172 -2799 -138
rect -2731 -172 -2715 -138
rect -2657 -172 -2641 -138
rect -2573 -172 -2557 -138
rect -2499 -172 -2483 -138
rect -2415 -172 -2399 -138
rect -2341 -172 -2325 -138
rect -2257 -172 -2241 -138
rect -2183 -172 -2167 -138
rect -2099 -172 -2083 -138
rect -2025 -172 -2009 -138
rect -1941 -172 -1925 -138
rect -1867 -172 -1851 -138
rect -1783 -172 -1767 -138
rect -1709 -172 -1693 -138
rect -1625 -172 -1609 -138
rect -1551 -172 -1535 -138
rect -1467 -172 -1451 -138
rect -1393 -172 -1377 -138
rect -1309 -172 -1293 -138
rect -1235 -172 -1219 -138
rect -1151 -172 -1135 -138
rect -1077 -172 -1061 -138
rect -993 -172 -977 -138
rect -919 -172 -903 -138
rect -835 -172 -819 -138
rect -761 -172 -745 -138
rect -677 -172 -661 -138
rect -603 -172 -587 -138
rect -519 -172 -503 -138
rect -445 -172 -429 -138
rect -361 -172 -345 -138
rect -287 -172 -271 -138
rect -203 -172 -187 -138
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 113 -172 129 -138
rect 187 -172 203 -138
rect 271 -172 287 -138
rect 345 -172 361 -138
rect 429 -172 445 -138
rect 503 -172 519 -138
rect 587 -172 603 -138
rect 661 -172 677 -138
rect 745 -172 761 -138
rect 819 -172 835 -138
rect 903 -172 919 -138
rect 977 -172 993 -138
rect 1061 -172 1077 -138
rect 1135 -172 1151 -138
rect 1219 -172 1235 -138
rect 1293 -172 1309 -138
rect 1377 -172 1393 -138
rect 1451 -172 1467 -138
rect 1535 -172 1551 -138
rect 1609 -172 1625 -138
rect 1693 -172 1709 -138
rect 1767 -172 1783 -138
rect 1851 -172 1867 -138
rect 1925 -172 1941 -138
rect 2009 -172 2025 -138
rect 2083 -172 2099 -138
rect 2167 -172 2183 -138
rect 2241 -172 2257 -138
rect 2325 -172 2341 -138
rect 2399 -172 2415 -138
rect 2483 -172 2499 -138
rect 2557 -172 2573 -138
rect 2641 -172 2657 -138
rect 2715 -172 2731 -138
rect 2799 -172 2815 -138
rect 2873 -172 2889 -138
rect 2957 -172 2973 -138
rect 3031 -172 3047 -138
rect 3115 -172 3131 -138
rect -3131 -280 -3115 -246
rect -3047 -280 -3031 -246
rect -2973 -280 -2957 -246
rect -2889 -280 -2873 -246
rect -2815 -280 -2799 -246
rect -2731 -280 -2715 -246
rect -2657 -280 -2641 -246
rect -2573 -280 -2557 -246
rect -2499 -280 -2483 -246
rect -2415 -280 -2399 -246
rect -2341 -280 -2325 -246
rect -2257 -280 -2241 -246
rect -2183 -280 -2167 -246
rect -2099 -280 -2083 -246
rect -2025 -280 -2009 -246
rect -1941 -280 -1925 -246
rect -1867 -280 -1851 -246
rect -1783 -280 -1767 -246
rect -1709 -280 -1693 -246
rect -1625 -280 -1609 -246
rect -1551 -280 -1535 -246
rect -1467 -280 -1451 -246
rect -1393 -280 -1377 -246
rect -1309 -280 -1293 -246
rect -1235 -280 -1219 -246
rect -1151 -280 -1135 -246
rect -1077 -280 -1061 -246
rect -993 -280 -977 -246
rect -919 -280 -903 -246
rect -835 -280 -819 -246
rect -761 -280 -745 -246
rect -677 -280 -661 -246
rect -603 -280 -587 -246
rect -519 -280 -503 -246
rect -445 -280 -429 -246
rect -361 -280 -345 -246
rect -287 -280 -271 -246
rect -203 -280 -187 -246
rect -129 -280 -113 -246
rect -45 -280 -29 -246
rect 29 -280 45 -246
rect 113 -280 129 -246
rect 187 -280 203 -246
rect 271 -280 287 -246
rect 345 -280 361 -246
rect 429 -280 445 -246
rect 503 -280 519 -246
rect 587 -280 603 -246
rect 661 -280 677 -246
rect 745 -280 761 -246
rect 819 -280 835 -246
rect 903 -280 919 -246
rect 977 -280 993 -246
rect 1061 -280 1077 -246
rect 1135 -280 1151 -246
rect 1219 -280 1235 -246
rect 1293 -280 1309 -246
rect 1377 -280 1393 -246
rect 1451 -280 1467 -246
rect 1535 -280 1551 -246
rect 1609 -280 1625 -246
rect 1693 -280 1709 -246
rect 1767 -280 1783 -246
rect 1851 -280 1867 -246
rect 1925 -280 1941 -246
rect 2009 -280 2025 -246
rect 2083 -280 2099 -246
rect 2167 -280 2183 -246
rect 2241 -280 2257 -246
rect 2325 -280 2341 -246
rect 2399 -280 2415 -246
rect 2483 -280 2499 -246
rect 2557 -280 2573 -246
rect 2641 -280 2657 -246
rect 2715 -280 2731 -246
rect 2799 -280 2815 -246
rect 2873 -280 2889 -246
rect 2957 -280 2973 -246
rect 3031 -280 3047 -246
rect 3115 -280 3131 -246
rect -3177 -330 -3143 -314
rect -3177 -522 -3143 -506
rect -3019 -330 -2985 -314
rect -3019 -522 -2985 -506
rect -2861 -330 -2827 -314
rect -2861 -522 -2827 -506
rect -2703 -330 -2669 -314
rect -2703 -522 -2669 -506
rect -2545 -330 -2511 -314
rect -2545 -522 -2511 -506
rect -2387 -330 -2353 -314
rect -2387 -522 -2353 -506
rect -2229 -330 -2195 -314
rect -2229 -522 -2195 -506
rect -2071 -330 -2037 -314
rect -2071 -522 -2037 -506
rect -1913 -330 -1879 -314
rect -1913 -522 -1879 -506
rect -1755 -330 -1721 -314
rect -1755 -522 -1721 -506
rect -1597 -330 -1563 -314
rect -1597 -522 -1563 -506
rect -1439 -330 -1405 -314
rect -1439 -522 -1405 -506
rect -1281 -330 -1247 -314
rect -1281 -522 -1247 -506
rect -1123 -330 -1089 -314
rect -1123 -522 -1089 -506
rect -965 -330 -931 -314
rect -965 -522 -931 -506
rect -807 -330 -773 -314
rect -807 -522 -773 -506
rect -649 -330 -615 -314
rect -649 -522 -615 -506
rect -491 -330 -457 -314
rect -491 -522 -457 -506
rect -333 -330 -299 -314
rect -333 -522 -299 -506
rect -175 -330 -141 -314
rect -175 -522 -141 -506
rect -17 -330 17 -314
rect -17 -522 17 -506
rect 141 -330 175 -314
rect 141 -522 175 -506
rect 299 -330 333 -314
rect 299 -522 333 -506
rect 457 -330 491 -314
rect 457 -522 491 -506
rect 615 -330 649 -314
rect 615 -522 649 -506
rect 773 -330 807 -314
rect 773 -522 807 -506
rect 931 -330 965 -314
rect 931 -522 965 -506
rect 1089 -330 1123 -314
rect 1089 -522 1123 -506
rect 1247 -330 1281 -314
rect 1247 -522 1281 -506
rect 1405 -330 1439 -314
rect 1405 -522 1439 -506
rect 1563 -330 1597 -314
rect 1563 -522 1597 -506
rect 1721 -330 1755 -314
rect 1721 -522 1755 -506
rect 1879 -330 1913 -314
rect 1879 -522 1913 -506
rect 2037 -330 2071 -314
rect 2037 -522 2071 -506
rect 2195 -330 2229 -314
rect 2195 -522 2229 -506
rect 2353 -330 2387 -314
rect 2353 -522 2387 -506
rect 2511 -330 2545 -314
rect 2511 -522 2545 -506
rect 2669 -330 2703 -314
rect 2669 -522 2703 -506
rect 2827 -330 2861 -314
rect 2827 -522 2861 -506
rect 2985 -330 3019 -314
rect 2985 -522 3019 -506
rect 3143 -330 3177 -314
rect 3143 -522 3177 -506
rect -3131 -590 -3115 -556
rect -3047 -590 -3031 -556
rect -2973 -590 -2957 -556
rect -2889 -590 -2873 -556
rect -2815 -590 -2799 -556
rect -2731 -590 -2715 -556
rect -2657 -590 -2641 -556
rect -2573 -590 -2557 -556
rect -2499 -590 -2483 -556
rect -2415 -590 -2399 -556
rect -2341 -590 -2325 -556
rect -2257 -590 -2241 -556
rect -2183 -590 -2167 -556
rect -2099 -590 -2083 -556
rect -2025 -590 -2009 -556
rect -1941 -590 -1925 -556
rect -1867 -590 -1851 -556
rect -1783 -590 -1767 -556
rect -1709 -590 -1693 -556
rect -1625 -590 -1609 -556
rect -1551 -590 -1535 -556
rect -1467 -590 -1451 -556
rect -1393 -590 -1377 -556
rect -1309 -590 -1293 -556
rect -1235 -590 -1219 -556
rect -1151 -590 -1135 -556
rect -1077 -590 -1061 -556
rect -993 -590 -977 -556
rect -919 -590 -903 -556
rect -835 -590 -819 -556
rect -761 -590 -745 -556
rect -677 -590 -661 -556
rect -603 -590 -587 -556
rect -519 -590 -503 -556
rect -445 -590 -429 -556
rect -361 -590 -345 -556
rect -287 -590 -271 -556
rect -203 -590 -187 -556
rect -129 -590 -113 -556
rect -45 -590 -29 -556
rect 29 -590 45 -556
rect 113 -590 129 -556
rect 187 -590 203 -556
rect 271 -590 287 -556
rect 345 -590 361 -556
rect 429 -590 445 -556
rect 503 -590 519 -556
rect 587 -590 603 -556
rect 661 -590 677 -556
rect 745 -590 761 -556
rect 819 -590 835 -556
rect 903 -590 919 -556
rect 977 -590 993 -556
rect 1061 -590 1077 -556
rect 1135 -590 1151 -556
rect 1219 -590 1235 -556
rect 1293 -590 1309 -556
rect 1377 -590 1393 -556
rect 1451 -590 1467 -556
rect 1535 -590 1551 -556
rect 1609 -590 1625 -556
rect 1693 -590 1709 -556
rect 1767 -590 1783 -556
rect 1851 -590 1867 -556
rect 1925 -590 1941 -556
rect 2009 -590 2025 -556
rect 2083 -590 2099 -556
rect 2167 -590 2183 -556
rect 2241 -590 2257 -556
rect 2325 -590 2341 -556
rect 2399 -590 2415 -556
rect 2483 -590 2499 -556
rect 2557 -590 2573 -556
rect 2641 -590 2657 -556
rect 2715 -590 2731 -556
rect 2799 -590 2815 -556
rect 2873 -590 2889 -556
rect 2957 -590 2973 -556
rect 3031 -590 3047 -556
rect 3115 -590 3131 -556
rect -3311 -694 -3277 -632
rect 3277 -694 3311 -632
rect -3311 -728 -3215 -694
rect 3215 -728 3311 -694
<< viali >>
rect -3115 556 -3047 590
rect -2957 556 -2889 590
rect -2799 556 -2731 590
rect -2641 556 -2573 590
rect -2483 556 -2415 590
rect -2325 556 -2257 590
rect -2167 556 -2099 590
rect -2009 556 -1941 590
rect -1851 556 -1783 590
rect -1693 556 -1625 590
rect -1535 556 -1467 590
rect -1377 556 -1309 590
rect -1219 556 -1151 590
rect -1061 556 -993 590
rect -903 556 -835 590
rect -745 556 -677 590
rect -587 556 -519 590
rect -429 556 -361 590
rect -271 556 -203 590
rect -113 556 -45 590
rect 45 556 113 590
rect 203 556 271 590
rect 361 556 429 590
rect 519 556 587 590
rect 677 556 745 590
rect 835 556 903 590
rect 993 556 1061 590
rect 1151 556 1219 590
rect 1309 556 1377 590
rect 1467 556 1535 590
rect 1625 556 1693 590
rect 1783 556 1851 590
rect 1941 556 2009 590
rect 2099 556 2167 590
rect 2257 556 2325 590
rect 2415 556 2483 590
rect 2573 556 2641 590
rect 2731 556 2799 590
rect 2889 556 2957 590
rect 3047 556 3115 590
rect -3177 330 -3143 506
rect -3019 330 -2985 506
rect -2861 330 -2827 506
rect -2703 330 -2669 506
rect -2545 330 -2511 506
rect -2387 330 -2353 506
rect -2229 330 -2195 506
rect -2071 330 -2037 506
rect -1913 330 -1879 506
rect -1755 330 -1721 506
rect -1597 330 -1563 506
rect -1439 330 -1405 506
rect -1281 330 -1247 506
rect -1123 330 -1089 506
rect -965 330 -931 506
rect -807 330 -773 506
rect -649 330 -615 506
rect -491 330 -457 506
rect -333 330 -299 506
rect -175 330 -141 506
rect -17 330 17 506
rect 141 330 175 506
rect 299 330 333 506
rect 457 330 491 506
rect 615 330 649 506
rect 773 330 807 506
rect 931 330 965 506
rect 1089 330 1123 506
rect 1247 330 1281 506
rect 1405 330 1439 506
rect 1563 330 1597 506
rect 1721 330 1755 506
rect 1879 330 1913 506
rect 2037 330 2071 506
rect 2195 330 2229 506
rect 2353 330 2387 506
rect 2511 330 2545 506
rect 2669 330 2703 506
rect 2827 330 2861 506
rect 2985 330 3019 506
rect 3143 330 3177 506
rect -3115 246 -3047 280
rect -2957 246 -2889 280
rect -2799 246 -2731 280
rect -2641 246 -2573 280
rect -2483 246 -2415 280
rect -2325 246 -2257 280
rect -2167 246 -2099 280
rect -2009 246 -1941 280
rect -1851 246 -1783 280
rect -1693 246 -1625 280
rect -1535 246 -1467 280
rect -1377 246 -1309 280
rect -1219 246 -1151 280
rect -1061 246 -993 280
rect -903 246 -835 280
rect -745 246 -677 280
rect -587 246 -519 280
rect -429 246 -361 280
rect -271 246 -203 280
rect -113 246 -45 280
rect 45 246 113 280
rect 203 246 271 280
rect 361 246 429 280
rect 519 246 587 280
rect 677 246 745 280
rect 835 246 903 280
rect 993 246 1061 280
rect 1151 246 1219 280
rect 1309 246 1377 280
rect 1467 246 1535 280
rect 1625 246 1693 280
rect 1783 246 1851 280
rect 1941 246 2009 280
rect 2099 246 2167 280
rect 2257 246 2325 280
rect 2415 246 2483 280
rect 2573 246 2641 280
rect 2731 246 2799 280
rect 2889 246 2957 280
rect 3047 246 3115 280
rect -3115 138 -3047 172
rect -2957 138 -2889 172
rect -2799 138 -2731 172
rect -2641 138 -2573 172
rect -2483 138 -2415 172
rect -2325 138 -2257 172
rect -2167 138 -2099 172
rect -2009 138 -1941 172
rect -1851 138 -1783 172
rect -1693 138 -1625 172
rect -1535 138 -1467 172
rect -1377 138 -1309 172
rect -1219 138 -1151 172
rect -1061 138 -993 172
rect -903 138 -835 172
rect -745 138 -677 172
rect -587 138 -519 172
rect -429 138 -361 172
rect -271 138 -203 172
rect -113 138 -45 172
rect 45 138 113 172
rect 203 138 271 172
rect 361 138 429 172
rect 519 138 587 172
rect 677 138 745 172
rect 835 138 903 172
rect 993 138 1061 172
rect 1151 138 1219 172
rect 1309 138 1377 172
rect 1467 138 1535 172
rect 1625 138 1693 172
rect 1783 138 1851 172
rect 1941 138 2009 172
rect 2099 138 2167 172
rect 2257 138 2325 172
rect 2415 138 2483 172
rect 2573 138 2641 172
rect 2731 138 2799 172
rect 2889 138 2957 172
rect 3047 138 3115 172
rect -3177 -88 -3143 88
rect -3019 -88 -2985 88
rect -2861 -88 -2827 88
rect -2703 -88 -2669 88
rect -2545 -88 -2511 88
rect -2387 -88 -2353 88
rect -2229 -88 -2195 88
rect -2071 -88 -2037 88
rect -1913 -88 -1879 88
rect -1755 -88 -1721 88
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
rect 1721 -88 1755 88
rect 1879 -88 1913 88
rect 2037 -88 2071 88
rect 2195 -88 2229 88
rect 2353 -88 2387 88
rect 2511 -88 2545 88
rect 2669 -88 2703 88
rect 2827 -88 2861 88
rect 2985 -88 3019 88
rect 3143 -88 3177 88
rect -3115 -172 -3047 -138
rect -2957 -172 -2889 -138
rect -2799 -172 -2731 -138
rect -2641 -172 -2573 -138
rect -2483 -172 -2415 -138
rect -2325 -172 -2257 -138
rect -2167 -172 -2099 -138
rect -2009 -172 -1941 -138
rect -1851 -172 -1783 -138
rect -1693 -172 -1625 -138
rect -1535 -172 -1467 -138
rect -1377 -172 -1309 -138
rect -1219 -172 -1151 -138
rect -1061 -172 -993 -138
rect -903 -172 -835 -138
rect -745 -172 -677 -138
rect -587 -172 -519 -138
rect -429 -172 -361 -138
rect -271 -172 -203 -138
rect -113 -172 -45 -138
rect 45 -172 113 -138
rect 203 -172 271 -138
rect 361 -172 429 -138
rect 519 -172 587 -138
rect 677 -172 745 -138
rect 835 -172 903 -138
rect 993 -172 1061 -138
rect 1151 -172 1219 -138
rect 1309 -172 1377 -138
rect 1467 -172 1535 -138
rect 1625 -172 1693 -138
rect 1783 -172 1851 -138
rect 1941 -172 2009 -138
rect 2099 -172 2167 -138
rect 2257 -172 2325 -138
rect 2415 -172 2483 -138
rect 2573 -172 2641 -138
rect 2731 -172 2799 -138
rect 2889 -172 2957 -138
rect 3047 -172 3115 -138
rect -3115 -280 -3047 -246
rect -2957 -280 -2889 -246
rect -2799 -280 -2731 -246
rect -2641 -280 -2573 -246
rect -2483 -280 -2415 -246
rect -2325 -280 -2257 -246
rect -2167 -280 -2099 -246
rect -2009 -280 -1941 -246
rect -1851 -280 -1783 -246
rect -1693 -280 -1625 -246
rect -1535 -280 -1467 -246
rect -1377 -280 -1309 -246
rect -1219 -280 -1151 -246
rect -1061 -280 -993 -246
rect -903 -280 -835 -246
rect -745 -280 -677 -246
rect -587 -280 -519 -246
rect -429 -280 -361 -246
rect -271 -280 -203 -246
rect -113 -280 -45 -246
rect 45 -280 113 -246
rect 203 -280 271 -246
rect 361 -280 429 -246
rect 519 -280 587 -246
rect 677 -280 745 -246
rect 835 -280 903 -246
rect 993 -280 1061 -246
rect 1151 -280 1219 -246
rect 1309 -280 1377 -246
rect 1467 -280 1535 -246
rect 1625 -280 1693 -246
rect 1783 -280 1851 -246
rect 1941 -280 2009 -246
rect 2099 -280 2167 -246
rect 2257 -280 2325 -246
rect 2415 -280 2483 -246
rect 2573 -280 2641 -246
rect 2731 -280 2799 -246
rect 2889 -280 2957 -246
rect 3047 -280 3115 -246
rect -3177 -506 -3143 -330
rect -3019 -506 -2985 -330
rect -2861 -506 -2827 -330
rect -2703 -506 -2669 -330
rect -2545 -506 -2511 -330
rect -2387 -506 -2353 -330
rect -2229 -506 -2195 -330
rect -2071 -506 -2037 -330
rect -1913 -506 -1879 -330
rect -1755 -506 -1721 -330
rect -1597 -506 -1563 -330
rect -1439 -506 -1405 -330
rect -1281 -506 -1247 -330
rect -1123 -506 -1089 -330
rect -965 -506 -931 -330
rect -807 -506 -773 -330
rect -649 -506 -615 -330
rect -491 -506 -457 -330
rect -333 -506 -299 -330
rect -175 -506 -141 -330
rect -17 -506 17 -330
rect 141 -506 175 -330
rect 299 -506 333 -330
rect 457 -506 491 -330
rect 615 -506 649 -330
rect 773 -506 807 -330
rect 931 -506 965 -330
rect 1089 -506 1123 -330
rect 1247 -506 1281 -330
rect 1405 -506 1439 -330
rect 1563 -506 1597 -330
rect 1721 -506 1755 -330
rect 1879 -506 1913 -330
rect 2037 -506 2071 -330
rect 2195 -506 2229 -330
rect 2353 -506 2387 -330
rect 2511 -506 2545 -330
rect 2669 -506 2703 -330
rect 2827 -506 2861 -330
rect 2985 -506 3019 -330
rect 3143 -506 3177 -330
rect -3115 -590 -3047 -556
rect -2957 -590 -2889 -556
rect -2799 -590 -2731 -556
rect -2641 -590 -2573 -556
rect -2483 -590 -2415 -556
rect -2325 -590 -2257 -556
rect -2167 -590 -2099 -556
rect -2009 -590 -1941 -556
rect -1851 -590 -1783 -556
rect -1693 -590 -1625 -556
rect -1535 -590 -1467 -556
rect -1377 -590 -1309 -556
rect -1219 -590 -1151 -556
rect -1061 -590 -993 -556
rect -903 -590 -835 -556
rect -745 -590 -677 -556
rect -587 -590 -519 -556
rect -429 -590 -361 -556
rect -271 -590 -203 -556
rect -113 -590 -45 -556
rect 45 -590 113 -556
rect 203 -590 271 -556
rect 361 -590 429 -556
rect 519 -590 587 -556
rect 677 -590 745 -556
rect 835 -590 903 -556
rect 993 -590 1061 -556
rect 1151 -590 1219 -556
rect 1309 -590 1377 -556
rect 1467 -590 1535 -556
rect 1625 -590 1693 -556
rect 1783 -590 1851 -556
rect 1941 -590 2009 -556
rect 2099 -590 2167 -556
rect 2257 -590 2325 -556
rect 2415 -590 2483 -556
rect 2573 -590 2641 -556
rect 2731 -590 2799 -556
rect 2889 -590 2957 -556
rect 3047 -590 3115 -556
<< metal1 >>
rect -3127 590 -3035 596
rect -3127 556 -3115 590
rect -3047 556 -3035 590
rect -3127 550 -3035 556
rect -2969 590 -2877 596
rect -2969 556 -2957 590
rect -2889 556 -2877 590
rect -2969 550 -2877 556
rect -2811 590 -2719 596
rect -2811 556 -2799 590
rect -2731 556 -2719 590
rect -2811 550 -2719 556
rect -2653 590 -2561 596
rect -2653 556 -2641 590
rect -2573 556 -2561 590
rect -2653 550 -2561 556
rect -2495 590 -2403 596
rect -2495 556 -2483 590
rect -2415 556 -2403 590
rect -2495 550 -2403 556
rect -2337 590 -2245 596
rect -2337 556 -2325 590
rect -2257 556 -2245 590
rect -2337 550 -2245 556
rect -2179 590 -2087 596
rect -2179 556 -2167 590
rect -2099 556 -2087 590
rect -2179 550 -2087 556
rect -2021 590 -1929 596
rect -2021 556 -2009 590
rect -1941 556 -1929 590
rect -2021 550 -1929 556
rect -1863 590 -1771 596
rect -1863 556 -1851 590
rect -1783 556 -1771 590
rect -1863 550 -1771 556
rect -1705 590 -1613 596
rect -1705 556 -1693 590
rect -1625 556 -1613 590
rect -1705 550 -1613 556
rect -1547 590 -1455 596
rect -1547 556 -1535 590
rect -1467 556 -1455 590
rect -1547 550 -1455 556
rect -1389 590 -1297 596
rect -1389 556 -1377 590
rect -1309 556 -1297 590
rect -1389 550 -1297 556
rect -1231 590 -1139 596
rect -1231 556 -1219 590
rect -1151 556 -1139 590
rect -1231 550 -1139 556
rect -1073 590 -981 596
rect -1073 556 -1061 590
rect -993 556 -981 590
rect -1073 550 -981 556
rect -915 590 -823 596
rect -915 556 -903 590
rect -835 556 -823 590
rect -915 550 -823 556
rect -757 590 -665 596
rect -757 556 -745 590
rect -677 556 -665 590
rect -757 550 -665 556
rect -599 590 -507 596
rect -599 556 -587 590
rect -519 556 -507 590
rect -599 550 -507 556
rect -441 590 -349 596
rect -441 556 -429 590
rect -361 556 -349 590
rect -441 550 -349 556
rect -283 590 -191 596
rect -283 556 -271 590
rect -203 556 -191 590
rect -283 550 -191 556
rect -125 590 -33 596
rect -125 556 -113 590
rect -45 556 -33 590
rect -125 550 -33 556
rect 33 590 125 596
rect 33 556 45 590
rect 113 556 125 590
rect 33 550 125 556
rect 191 590 283 596
rect 191 556 203 590
rect 271 556 283 590
rect 191 550 283 556
rect 349 590 441 596
rect 349 556 361 590
rect 429 556 441 590
rect 349 550 441 556
rect 507 590 599 596
rect 507 556 519 590
rect 587 556 599 590
rect 507 550 599 556
rect 665 590 757 596
rect 665 556 677 590
rect 745 556 757 590
rect 665 550 757 556
rect 823 590 915 596
rect 823 556 835 590
rect 903 556 915 590
rect 823 550 915 556
rect 981 590 1073 596
rect 981 556 993 590
rect 1061 556 1073 590
rect 981 550 1073 556
rect 1139 590 1231 596
rect 1139 556 1151 590
rect 1219 556 1231 590
rect 1139 550 1231 556
rect 1297 590 1389 596
rect 1297 556 1309 590
rect 1377 556 1389 590
rect 1297 550 1389 556
rect 1455 590 1547 596
rect 1455 556 1467 590
rect 1535 556 1547 590
rect 1455 550 1547 556
rect 1613 590 1705 596
rect 1613 556 1625 590
rect 1693 556 1705 590
rect 1613 550 1705 556
rect 1771 590 1863 596
rect 1771 556 1783 590
rect 1851 556 1863 590
rect 1771 550 1863 556
rect 1929 590 2021 596
rect 1929 556 1941 590
rect 2009 556 2021 590
rect 1929 550 2021 556
rect 2087 590 2179 596
rect 2087 556 2099 590
rect 2167 556 2179 590
rect 2087 550 2179 556
rect 2245 590 2337 596
rect 2245 556 2257 590
rect 2325 556 2337 590
rect 2245 550 2337 556
rect 2403 590 2495 596
rect 2403 556 2415 590
rect 2483 556 2495 590
rect 2403 550 2495 556
rect 2561 590 2653 596
rect 2561 556 2573 590
rect 2641 556 2653 590
rect 2561 550 2653 556
rect 2719 590 2811 596
rect 2719 556 2731 590
rect 2799 556 2811 590
rect 2719 550 2811 556
rect 2877 590 2969 596
rect 2877 556 2889 590
rect 2957 556 2969 590
rect 2877 550 2969 556
rect 3035 590 3127 596
rect 3035 556 3047 590
rect 3115 556 3127 590
rect 3035 550 3127 556
rect -3183 506 -3137 518
rect -3183 330 -3177 506
rect -3143 330 -3137 506
rect -3183 318 -3137 330
rect -3025 506 -2979 518
rect -3025 330 -3019 506
rect -2985 330 -2979 506
rect -3025 318 -2979 330
rect -2867 506 -2821 518
rect -2867 330 -2861 506
rect -2827 330 -2821 506
rect -2867 318 -2821 330
rect -2709 506 -2663 518
rect -2709 330 -2703 506
rect -2669 330 -2663 506
rect -2709 318 -2663 330
rect -2551 506 -2505 518
rect -2551 330 -2545 506
rect -2511 330 -2505 506
rect -2551 318 -2505 330
rect -2393 506 -2347 518
rect -2393 330 -2387 506
rect -2353 330 -2347 506
rect -2393 318 -2347 330
rect -2235 506 -2189 518
rect -2235 330 -2229 506
rect -2195 330 -2189 506
rect -2235 318 -2189 330
rect -2077 506 -2031 518
rect -2077 330 -2071 506
rect -2037 330 -2031 506
rect -2077 318 -2031 330
rect -1919 506 -1873 518
rect -1919 330 -1913 506
rect -1879 330 -1873 506
rect -1919 318 -1873 330
rect -1761 506 -1715 518
rect -1761 330 -1755 506
rect -1721 330 -1715 506
rect -1761 318 -1715 330
rect -1603 506 -1557 518
rect -1603 330 -1597 506
rect -1563 330 -1557 506
rect -1603 318 -1557 330
rect -1445 506 -1399 518
rect -1445 330 -1439 506
rect -1405 330 -1399 506
rect -1445 318 -1399 330
rect -1287 506 -1241 518
rect -1287 330 -1281 506
rect -1247 330 -1241 506
rect -1287 318 -1241 330
rect -1129 506 -1083 518
rect -1129 330 -1123 506
rect -1089 330 -1083 506
rect -1129 318 -1083 330
rect -971 506 -925 518
rect -971 330 -965 506
rect -931 330 -925 506
rect -971 318 -925 330
rect -813 506 -767 518
rect -813 330 -807 506
rect -773 330 -767 506
rect -813 318 -767 330
rect -655 506 -609 518
rect -655 330 -649 506
rect -615 330 -609 506
rect -655 318 -609 330
rect -497 506 -451 518
rect -497 330 -491 506
rect -457 330 -451 506
rect -497 318 -451 330
rect -339 506 -293 518
rect -339 330 -333 506
rect -299 330 -293 506
rect -339 318 -293 330
rect -181 506 -135 518
rect -181 330 -175 506
rect -141 330 -135 506
rect -181 318 -135 330
rect -23 506 23 518
rect -23 330 -17 506
rect 17 330 23 506
rect -23 318 23 330
rect 135 506 181 518
rect 135 330 141 506
rect 175 330 181 506
rect 135 318 181 330
rect 293 506 339 518
rect 293 330 299 506
rect 333 330 339 506
rect 293 318 339 330
rect 451 506 497 518
rect 451 330 457 506
rect 491 330 497 506
rect 451 318 497 330
rect 609 506 655 518
rect 609 330 615 506
rect 649 330 655 506
rect 609 318 655 330
rect 767 506 813 518
rect 767 330 773 506
rect 807 330 813 506
rect 767 318 813 330
rect 925 506 971 518
rect 925 330 931 506
rect 965 330 971 506
rect 925 318 971 330
rect 1083 506 1129 518
rect 1083 330 1089 506
rect 1123 330 1129 506
rect 1083 318 1129 330
rect 1241 506 1287 518
rect 1241 330 1247 506
rect 1281 330 1287 506
rect 1241 318 1287 330
rect 1399 506 1445 518
rect 1399 330 1405 506
rect 1439 330 1445 506
rect 1399 318 1445 330
rect 1557 506 1603 518
rect 1557 330 1563 506
rect 1597 330 1603 506
rect 1557 318 1603 330
rect 1715 506 1761 518
rect 1715 330 1721 506
rect 1755 330 1761 506
rect 1715 318 1761 330
rect 1873 506 1919 518
rect 1873 330 1879 506
rect 1913 330 1919 506
rect 1873 318 1919 330
rect 2031 506 2077 518
rect 2031 330 2037 506
rect 2071 330 2077 506
rect 2031 318 2077 330
rect 2189 506 2235 518
rect 2189 330 2195 506
rect 2229 330 2235 506
rect 2189 318 2235 330
rect 2347 506 2393 518
rect 2347 330 2353 506
rect 2387 330 2393 506
rect 2347 318 2393 330
rect 2505 506 2551 518
rect 2505 330 2511 506
rect 2545 330 2551 506
rect 2505 318 2551 330
rect 2663 506 2709 518
rect 2663 330 2669 506
rect 2703 330 2709 506
rect 2663 318 2709 330
rect 2821 506 2867 518
rect 2821 330 2827 506
rect 2861 330 2867 506
rect 2821 318 2867 330
rect 2979 506 3025 518
rect 2979 330 2985 506
rect 3019 330 3025 506
rect 2979 318 3025 330
rect 3137 506 3183 518
rect 3137 330 3143 506
rect 3177 330 3183 506
rect 3137 318 3183 330
rect -3127 280 -3035 286
rect -3127 246 -3115 280
rect -3047 246 -3035 280
rect -3127 240 -3035 246
rect -2969 280 -2877 286
rect -2969 246 -2957 280
rect -2889 246 -2877 280
rect -2969 240 -2877 246
rect -2811 280 -2719 286
rect -2811 246 -2799 280
rect -2731 246 -2719 280
rect -2811 240 -2719 246
rect -2653 280 -2561 286
rect -2653 246 -2641 280
rect -2573 246 -2561 280
rect -2653 240 -2561 246
rect -2495 280 -2403 286
rect -2495 246 -2483 280
rect -2415 246 -2403 280
rect -2495 240 -2403 246
rect -2337 280 -2245 286
rect -2337 246 -2325 280
rect -2257 246 -2245 280
rect -2337 240 -2245 246
rect -2179 280 -2087 286
rect -2179 246 -2167 280
rect -2099 246 -2087 280
rect -2179 240 -2087 246
rect -2021 280 -1929 286
rect -2021 246 -2009 280
rect -1941 246 -1929 280
rect -2021 240 -1929 246
rect -1863 280 -1771 286
rect -1863 246 -1851 280
rect -1783 246 -1771 280
rect -1863 240 -1771 246
rect -1705 280 -1613 286
rect -1705 246 -1693 280
rect -1625 246 -1613 280
rect -1705 240 -1613 246
rect -1547 280 -1455 286
rect -1547 246 -1535 280
rect -1467 246 -1455 280
rect -1547 240 -1455 246
rect -1389 280 -1297 286
rect -1389 246 -1377 280
rect -1309 246 -1297 280
rect -1389 240 -1297 246
rect -1231 280 -1139 286
rect -1231 246 -1219 280
rect -1151 246 -1139 280
rect -1231 240 -1139 246
rect -1073 280 -981 286
rect -1073 246 -1061 280
rect -993 246 -981 280
rect -1073 240 -981 246
rect -915 280 -823 286
rect -915 246 -903 280
rect -835 246 -823 280
rect -915 240 -823 246
rect -757 280 -665 286
rect -757 246 -745 280
rect -677 246 -665 280
rect -757 240 -665 246
rect -599 280 -507 286
rect -599 246 -587 280
rect -519 246 -507 280
rect -599 240 -507 246
rect -441 280 -349 286
rect -441 246 -429 280
rect -361 246 -349 280
rect -441 240 -349 246
rect -283 280 -191 286
rect -283 246 -271 280
rect -203 246 -191 280
rect -283 240 -191 246
rect -125 280 -33 286
rect -125 246 -113 280
rect -45 246 -33 280
rect -125 240 -33 246
rect 33 280 125 286
rect 33 246 45 280
rect 113 246 125 280
rect 33 240 125 246
rect 191 280 283 286
rect 191 246 203 280
rect 271 246 283 280
rect 191 240 283 246
rect 349 280 441 286
rect 349 246 361 280
rect 429 246 441 280
rect 349 240 441 246
rect 507 280 599 286
rect 507 246 519 280
rect 587 246 599 280
rect 507 240 599 246
rect 665 280 757 286
rect 665 246 677 280
rect 745 246 757 280
rect 665 240 757 246
rect 823 280 915 286
rect 823 246 835 280
rect 903 246 915 280
rect 823 240 915 246
rect 981 280 1073 286
rect 981 246 993 280
rect 1061 246 1073 280
rect 981 240 1073 246
rect 1139 280 1231 286
rect 1139 246 1151 280
rect 1219 246 1231 280
rect 1139 240 1231 246
rect 1297 280 1389 286
rect 1297 246 1309 280
rect 1377 246 1389 280
rect 1297 240 1389 246
rect 1455 280 1547 286
rect 1455 246 1467 280
rect 1535 246 1547 280
rect 1455 240 1547 246
rect 1613 280 1705 286
rect 1613 246 1625 280
rect 1693 246 1705 280
rect 1613 240 1705 246
rect 1771 280 1863 286
rect 1771 246 1783 280
rect 1851 246 1863 280
rect 1771 240 1863 246
rect 1929 280 2021 286
rect 1929 246 1941 280
rect 2009 246 2021 280
rect 1929 240 2021 246
rect 2087 280 2179 286
rect 2087 246 2099 280
rect 2167 246 2179 280
rect 2087 240 2179 246
rect 2245 280 2337 286
rect 2245 246 2257 280
rect 2325 246 2337 280
rect 2245 240 2337 246
rect 2403 280 2495 286
rect 2403 246 2415 280
rect 2483 246 2495 280
rect 2403 240 2495 246
rect 2561 280 2653 286
rect 2561 246 2573 280
rect 2641 246 2653 280
rect 2561 240 2653 246
rect 2719 280 2811 286
rect 2719 246 2731 280
rect 2799 246 2811 280
rect 2719 240 2811 246
rect 2877 280 2969 286
rect 2877 246 2889 280
rect 2957 246 2969 280
rect 2877 240 2969 246
rect 3035 280 3127 286
rect 3035 246 3047 280
rect 3115 246 3127 280
rect 3035 240 3127 246
rect -3127 172 -3035 178
rect -3127 138 -3115 172
rect -3047 138 -3035 172
rect -3127 132 -3035 138
rect -2969 172 -2877 178
rect -2969 138 -2957 172
rect -2889 138 -2877 172
rect -2969 132 -2877 138
rect -2811 172 -2719 178
rect -2811 138 -2799 172
rect -2731 138 -2719 172
rect -2811 132 -2719 138
rect -2653 172 -2561 178
rect -2653 138 -2641 172
rect -2573 138 -2561 172
rect -2653 132 -2561 138
rect -2495 172 -2403 178
rect -2495 138 -2483 172
rect -2415 138 -2403 172
rect -2495 132 -2403 138
rect -2337 172 -2245 178
rect -2337 138 -2325 172
rect -2257 138 -2245 172
rect -2337 132 -2245 138
rect -2179 172 -2087 178
rect -2179 138 -2167 172
rect -2099 138 -2087 172
rect -2179 132 -2087 138
rect -2021 172 -1929 178
rect -2021 138 -2009 172
rect -1941 138 -1929 172
rect -2021 132 -1929 138
rect -1863 172 -1771 178
rect -1863 138 -1851 172
rect -1783 138 -1771 172
rect -1863 132 -1771 138
rect -1705 172 -1613 178
rect -1705 138 -1693 172
rect -1625 138 -1613 172
rect -1705 132 -1613 138
rect -1547 172 -1455 178
rect -1547 138 -1535 172
rect -1467 138 -1455 172
rect -1547 132 -1455 138
rect -1389 172 -1297 178
rect -1389 138 -1377 172
rect -1309 138 -1297 172
rect -1389 132 -1297 138
rect -1231 172 -1139 178
rect -1231 138 -1219 172
rect -1151 138 -1139 172
rect -1231 132 -1139 138
rect -1073 172 -981 178
rect -1073 138 -1061 172
rect -993 138 -981 172
rect -1073 132 -981 138
rect -915 172 -823 178
rect -915 138 -903 172
rect -835 138 -823 172
rect -915 132 -823 138
rect -757 172 -665 178
rect -757 138 -745 172
rect -677 138 -665 172
rect -757 132 -665 138
rect -599 172 -507 178
rect -599 138 -587 172
rect -519 138 -507 172
rect -599 132 -507 138
rect -441 172 -349 178
rect -441 138 -429 172
rect -361 138 -349 172
rect -441 132 -349 138
rect -283 172 -191 178
rect -283 138 -271 172
rect -203 138 -191 172
rect -283 132 -191 138
rect -125 172 -33 178
rect -125 138 -113 172
rect -45 138 -33 172
rect -125 132 -33 138
rect 33 172 125 178
rect 33 138 45 172
rect 113 138 125 172
rect 33 132 125 138
rect 191 172 283 178
rect 191 138 203 172
rect 271 138 283 172
rect 191 132 283 138
rect 349 172 441 178
rect 349 138 361 172
rect 429 138 441 172
rect 349 132 441 138
rect 507 172 599 178
rect 507 138 519 172
rect 587 138 599 172
rect 507 132 599 138
rect 665 172 757 178
rect 665 138 677 172
rect 745 138 757 172
rect 665 132 757 138
rect 823 172 915 178
rect 823 138 835 172
rect 903 138 915 172
rect 823 132 915 138
rect 981 172 1073 178
rect 981 138 993 172
rect 1061 138 1073 172
rect 981 132 1073 138
rect 1139 172 1231 178
rect 1139 138 1151 172
rect 1219 138 1231 172
rect 1139 132 1231 138
rect 1297 172 1389 178
rect 1297 138 1309 172
rect 1377 138 1389 172
rect 1297 132 1389 138
rect 1455 172 1547 178
rect 1455 138 1467 172
rect 1535 138 1547 172
rect 1455 132 1547 138
rect 1613 172 1705 178
rect 1613 138 1625 172
rect 1693 138 1705 172
rect 1613 132 1705 138
rect 1771 172 1863 178
rect 1771 138 1783 172
rect 1851 138 1863 172
rect 1771 132 1863 138
rect 1929 172 2021 178
rect 1929 138 1941 172
rect 2009 138 2021 172
rect 1929 132 2021 138
rect 2087 172 2179 178
rect 2087 138 2099 172
rect 2167 138 2179 172
rect 2087 132 2179 138
rect 2245 172 2337 178
rect 2245 138 2257 172
rect 2325 138 2337 172
rect 2245 132 2337 138
rect 2403 172 2495 178
rect 2403 138 2415 172
rect 2483 138 2495 172
rect 2403 132 2495 138
rect 2561 172 2653 178
rect 2561 138 2573 172
rect 2641 138 2653 172
rect 2561 132 2653 138
rect 2719 172 2811 178
rect 2719 138 2731 172
rect 2799 138 2811 172
rect 2719 132 2811 138
rect 2877 172 2969 178
rect 2877 138 2889 172
rect 2957 138 2969 172
rect 2877 132 2969 138
rect 3035 172 3127 178
rect 3035 138 3047 172
rect 3115 138 3127 172
rect 3035 132 3127 138
rect -3183 88 -3137 100
rect -3183 -88 -3177 88
rect -3143 -88 -3137 88
rect -3183 -100 -3137 -88
rect -3025 88 -2979 100
rect -3025 -88 -3019 88
rect -2985 -88 -2979 88
rect -3025 -100 -2979 -88
rect -2867 88 -2821 100
rect -2867 -88 -2861 88
rect -2827 -88 -2821 88
rect -2867 -100 -2821 -88
rect -2709 88 -2663 100
rect -2709 -88 -2703 88
rect -2669 -88 -2663 88
rect -2709 -100 -2663 -88
rect -2551 88 -2505 100
rect -2551 -88 -2545 88
rect -2511 -88 -2505 88
rect -2551 -100 -2505 -88
rect -2393 88 -2347 100
rect -2393 -88 -2387 88
rect -2353 -88 -2347 88
rect -2393 -100 -2347 -88
rect -2235 88 -2189 100
rect -2235 -88 -2229 88
rect -2195 -88 -2189 88
rect -2235 -100 -2189 -88
rect -2077 88 -2031 100
rect -2077 -88 -2071 88
rect -2037 -88 -2031 88
rect -2077 -100 -2031 -88
rect -1919 88 -1873 100
rect -1919 -88 -1913 88
rect -1879 -88 -1873 88
rect -1919 -100 -1873 -88
rect -1761 88 -1715 100
rect -1761 -88 -1755 88
rect -1721 -88 -1715 88
rect -1761 -100 -1715 -88
rect -1603 88 -1557 100
rect -1603 -88 -1597 88
rect -1563 -88 -1557 88
rect -1603 -100 -1557 -88
rect -1445 88 -1399 100
rect -1445 -88 -1439 88
rect -1405 -88 -1399 88
rect -1445 -100 -1399 -88
rect -1287 88 -1241 100
rect -1287 -88 -1281 88
rect -1247 -88 -1241 88
rect -1287 -100 -1241 -88
rect -1129 88 -1083 100
rect -1129 -88 -1123 88
rect -1089 -88 -1083 88
rect -1129 -100 -1083 -88
rect -971 88 -925 100
rect -971 -88 -965 88
rect -931 -88 -925 88
rect -971 -100 -925 -88
rect -813 88 -767 100
rect -813 -88 -807 88
rect -773 -88 -767 88
rect -813 -100 -767 -88
rect -655 88 -609 100
rect -655 -88 -649 88
rect -615 -88 -609 88
rect -655 -100 -609 -88
rect -497 88 -451 100
rect -497 -88 -491 88
rect -457 -88 -451 88
rect -497 -100 -451 -88
rect -339 88 -293 100
rect -339 -88 -333 88
rect -299 -88 -293 88
rect -339 -100 -293 -88
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect 293 88 339 100
rect 293 -88 299 88
rect 333 -88 339 88
rect 293 -100 339 -88
rect 451 88 497 100
rect 451 -88 457 88
rect 491 -88 497 88
rect 451 -100 497 -88
rect 609 88 655 100
rect 609 -88 615 88
rect 649 -88 655 88
rect 609 -100 655 -88
rect 767 88 813 100
rect 767 -88 773 88
rect 807 -88 813 88
rect 767 -100 813 -88
rect 925 88 971 100
rect 925 -88 931 88
rect 965 -88 971 88
rect 925 -100 971 -88
rect 1083 88 1129 100
rect 1083 -88 1089 88
rect 1123 -88 1129 88
rect 1083 -100 1129 -88
rect 1241 88 1287 100
rect 1241 -88 1247 88
rect 1281 -88 1287 88
rect 1241 -100 1287 -88
rect 1399 88 1445 100
rect 1399 -88 1405 88
rect 1439 -88 1445 88
rect 1399 -100 1445 -88
rect 1557 88 1603 100
rect 1557 -88 1563 88
rect 1597 -88 1603 88
rect 1557 -100 1603 -88
rect 1715 88 1761 100
rect 1715 -88 1721 88
rect 1755 -88 1761 88
rect 1715 -100 1761 -88
rect 1873 88 1919 100
rect 1873 -88 1879 88
rect 1913 -88 1919 88
rect 1873 -100 1919 -88
rect 2031 88 2077 100
rect 2031 -88 2037 88
rect 2071 -88 2077 88
rect 2031 -100 2077 -88
rect 2189 88 2235 100
rect 2189 -88 2195 88
rect 2229 -88 2235 88
rect 2189 -100 2235 -88
rect 2347 88 2393 100
rect 2347 -88 2353 88
rect 2387 -88 2393 88
rect 2347 -100 2393 -88
rect 2505 88 2551 100
rect 2505 -88 2511 88
rect 2545 -88 2551 88
rect 2505 -100 2551 -88
rect 2663 88 2709 100
rect 2663 -88 2669 88
rect 2703 -88 2709 88
rect 2663 -100 2709 -88
rect 2821 88 2867 100
rect 2821 -88 2827 88
rect 2861 -88 2867 88
rect 2821 -100 2867 -88
rect 2979 88 3025 100
rect 2979 -88 2985 88
rect 3019 -88 3025 88
rect 2979 -100 3025 -88
rect 3137 88 3183 100
rect 3137 -88 3143 88
rect 3177 -88 3183 88
rect 3137 -100 3183 -88
rect -3127 -138 -3035 -132
rect -3127 -172 -3115 -138
rect -3047 -172 -3035 -138
rect -3127 -178 -3035 -172
rect -2969 -138 -2877 -132
rect -2969 -172 -2957 -138
rect -2889 -172 -2877 -138
rect -2969 -178 -2877 -172
rect -2811 -138 -2719 -132
rect -2811 -172 -2799 -138
rect -2731 -172 -2719 -138
rect -2811 -178 -2719 -172
rect -2653 -138 -2561 -132
rect -2653 -172 -2641 -138
rect -2573 -172 -2561 -138
rect -2653 -178 -2561 -172
rect -2495 -138 -2403 -132
rect -2495 -172 -2483 -138
rect -2415 -172 -2403 -138
rect -2495 -178 -2403 -172
rect -2337 -138 -2245 -132
rect -2337 -172 -2325 -138
rect -2257 -172 -2245 -138
rect -2337 -178 -2245 -172
rect -2179 -138 -2087 -132
rect -2179 -172 -2167 -138
rect -2099 -172 -2087 -138
rect -2179 -178 -2087 -172
rect -2021 -138 -1929 -132
rect -2021 -172 -2009 -138
rect -1941 -172 -1929 -138
rect -2021 -178 -1929 -172
rect -1863 -138 -1771 -132
rect -1863 -172 -1851 -138
rect -1783 -172 -1771 -138
rect -1863 -178 -1771 -172
rect -1705 -138 -1613 -132
rect -1705 -172 -1693 -138
rect -1625 -172 -1613 -138
rect -1705 -178 -1613 -172
rect -1547 -138 -1455 -132
rect -1547 -172 -1535 -138
rect -1467 -172 -1455 -138
rect -1547 -178 -1455 -172
rect -1389 -138 -1297 -132
rect -1389 -172 -1377 -138
rect -1309 -172 -1297 -138
rect -1389 -178 -1297 -172
rect -1231 -138 -1139 -132
rect -1231 -172 -1219 -138
rect -1151 -172 -1139 -138
rect -1231 -178 -1139 -172
rect -1073 -138 -981 -132
rect -1073 -172 -1061 -138
rect -993 -172 -981 -138
rect -1073 -178 -981 -172
rect -915 -138 -823 -132
rect -915 -172 -903 -138
rect -835 -172 -823 -138
rect -915 -178 -823 -172
rect -757 -138 -665 -132
rect -757 -172 -745 -138
rect -677 -172 -665 -138
rect -757 -178 -665 -172
rect -599 -138 -507 -132
rect -599 -172 -587 -138
rect -519 -172 -507 -138
rect -599 -178 -507 -172
rect -441 -138 -349 -132
rect -441 -172 -429 -138
rect -361 -172 -349 -138
rect -441 -178 -349 -172
rect -283 -138 -191 -132
rect -283 -172 -271 -138
rect -203 -172 -191 -138
rect -283 -178 -191 -172
rect -125 -138 -33 -132
rect -125 -172 -113 -138
rect -45 -172 -33 -138
rect -125 -178 -33 -172
rect 33 -138 125 -132
rect 33 -172 45 -138
rect 113 -172 125 -138
rect 33 -178 125 -172
rect 191 -138 283 -132
rect 191 -172 203 -138
rect 271 -172 283 -138
rect 191 -178 283 -172
rect 349 -138 441 -132
rect 349 -172 361 -138
rect 429 -172 441 -138
rect 349 -178 441 -172
rect 507 -138 599 -132
rect 507 -172 519 -138
rect 587 -172 599 -138
rect 507 -178 599 -172
rect 665 -138 757 -132
rect 665 -172 677 -138
rect 745 -172 757 -138
rect 665 -178 757 -172
rect 823 -138 915 -132
rect 823 -172 835 -138
rect 903 -172 915 -138
rect 823 -178 915 -172
rect 981 -138 1073 -132
rect 981 -172 993 -138
rect 1061 -172 1073 -138
rect 981 -178 1073 -172
rect 1139 -138 1231 -132
rect 1139 -172 1151 -138
rect 1219 -172 1231 -138
rect 1139 -178 1231 -172
rect 1297 -138 1389 -132
rect 1297 -172 1309 -138
rect 1377 -172 1389 -138
rect 1297 -178 1389 -172
rect 1455 -138 1547 -132
rect 1455 -172 1467 -138
rect 1535 -172 1547 -138
rect 1455 -178 1547 -172
rect 1613 -138 1705 -132
rect 1613 -172 1625 -138
rect 1693 -172 1705 -138
rect 1613 -178 1705 -172
rect 1771 -138 1863 -132
rect 1771 -172 1783 -138
rect 1851 -172 1863 -138
rect 1771 -178 1863 -172
rect 1929 -138 2021 -132
rect 1929 -172 1941 -138
rect 2009 -172 2021 -138
rect 1929 -178 2021 -172
rect 2087 -138 2179 -132
rect 2087 -172 2099 -138
rect 2167 -172 2179 -138
rect 2087 -178 2179 -172
rect 2245 -138 2337 -132
rect 2245 -172 2257 -138
rect 2325 -172 2337 -138
rect 2245 -178 2337 -172
rect 2403 -138 2495 -132
rect 2403 -172 2415 -138
rect 2483 -172 2495 -138
rect 2403 -178 2495 -172
rect 2561 -138 2653 -132
rect 2561 -172 2573 -138
rect 2641 -172 2653 -138
rect 2561 -178 2653 -172
rect 2719 -138 2811 -132
rect 2719 -172 2731 -138
rect 2799 -172 2811 -138
rect 2719 -178 2811 -172
rect 2877 -138 2969 -132
rect 2877 -172 2889 -138
rect 2957 -172 2969 -138
rect 2877 -178 2969 -172
rect 3035 -138 3127 -132
rect 3035 -172 3047 -138
rect 3115 -172 3127 -138
rect 3035 -178 3127 -172
rect -3127 -246 -3035 -240
rect -3127 -280 -3115 -246
rect -3047 -280 -3035 -246
rect -3127 -286 -3035 -280
rect -2969 -246 -2877 -240
rect -2969 -280 -2957 -246
rect -2889 -280 -2877 -246
rect -2969 -286 -2877 -280
rect -2811 -246 -2719 -240
rect -2811 -280 -2799 -246
rect -2731 -280 -2719 -246
rect -2811 -286 -2719 -280
rect -2653 -246 -2561 -240
rect -2653 -280 -2641 -246
rect -2573 -280 -2561 -246
rect -2653 -286 -2561 -280
rect -2495 -246 -2403 -240
rect -2495 -280 -2483 -246
rect -2415 -280 -2403 -246
rect -2495 -286 -2403 -280
rect -2337 -246 -2245 -240
rect -2337 -280 -2325 -246
rect -2257 -280 -2245 -246
rect -2337 -286 -2245 -280
rect -2179 -246 -2087 -240
rect -2179 -280 -2167 -246
rect -2099 -280 -2087 -246
rect -2179 -286 -2087 -280
rect -2021 -246 -1929 -240
rect -2021 -280 -2009 -246
rect -1941 -280 -1929 -246
rect -2021 -286 -1929 -280
rect -1863 -246 -1771 -240
rect -1863 -280 -1851 -246
rect -1783 -280 -1771 -246
rect -1863 -286 -1771 -280
rect -1705 -246 -1613 -240
rect -1705 -280 -1693 -246
rect -1625 -280 -1613 -246
rect -1705 -286 -1613 -280
rect -1547 -246 -1455 -240
rect -1547 -280 -1535 -246
rect -1467 -280 -1455 -246
rect -1547 -286 -1455 -280
rect -1389 -246 -1297 -240
rect -1389 -280 -1377 -246
rect -1309 -280 -1297 -246
rect -1389 -286 -1297 -280
rect -1231 -246 -1139 -240
rect -1231 -280 -1219 -246
rect -1151 -280 -1139 -246
rect -1231 -286 -1139 -280
rect -1073 -246 -981 -240
rect -1073 -280 -1061 -246
rect -993 -280 -981 -246
rect -1073 -286 -981 -280
rect -915 -246 -823 -240
rect -915 -280 -903 -246
rect -835 -280 -823 -246
rect -915 -286 -823 -280
rect -757 -246 -665 -240
rect -757 -280 -745 -246
rect -677 -280 -665 -246
rect -757 -286 -665 -280
rect -599 -246 -507 -240
rect -599 -280 -587 -246
rect -519 -280 -507 -246
rect -599 -286 -507 -280
rect -441 -246 -349 -240
rect -441 -280 -429 -246
rect -361 -280 -349 -246
rect -441 -286 -349 -280
rect -283 -246 -191 -240
rect -283 -280 -271 -246
rect -203 -280 -191 -246
rect -283 -286 -191 -280
rect -125 -246 -33 -240
rect -125 -280 -113 -246
rect -45 -280 -33 -246
rect -125 -286 -33 -280
rect 33 -246 125 -240
rect 33 -280 45 -246
rect 113 -280 125 -246
rect 33 -286 125 -280
rect 191 -246 283 -240
rect 191 -280 203 -246
rect 271 -280 283 -246
rect 191 -286 283 -280
rect 349 -246 441 -240
rect 349 -280 361 -246
rect 429 -280 441 -246
rect 349 -286 441 -280
rect 507 -246 599 -240
rect 507 -280 519 -246
rect 587 -280 599 -246
rect 507 -286 599 -280
rect 665 -246 757 -240
rect 665 -280 677 -246
rect 745 -280 757 -246
rect 665 -286 757 -280
rect 823 -246 915 -240
rect 823 -280 835 -246
rect 903 -280 915 -246
rect 823 -286 915 -280
rect 981 -246 1073 -240
rect 981 -280 993 -246
rect 1061 -280 1073 -246
rect 981 -286 1073 -280
rect 1139 -246 1231 -240
rect 1139 -280 1151 -246
rect 1219 -280 1231 -246
rect 1139 -286 1231 -280
rect 1297 -246 1389 -240
rect 1297 -280 1309 -246
rect 1377 -280 1389 -246
rect 1297 -286 1389 -280
rect 1455 -246 1547 -240
rect 1455 -280 1467 -246
rect 1535 -280 1547 -246
rect 1455 -286 1547 -280
rect 1613 -246 1705 -240
rect 1613 -280 1625 -246
rect 1693 -280 1705 -246
rect 1613 -286 1705 -280
rect 1771 -246 1863 -240
rect 1771 -280 1783 -246
rect 1851 -280 1863 -246
rect 1771 -286 1863 -280
rect 1929 -246 2021 -240
rect 1929 -280 1941 -246
rect 2009 -280 2021 -246
rect 1929 -286 2021 -280
rect 2087 -246 2179 -240
rect 2087 -280 2099 -246
rect 2167 -280 2179 -246
rect 2087 -286 2179 -280
rect 2245 -246 2337 -240
rect 2245 -280 2257 -246
rect 2325 -280 2337 -246
rect 2245 -286 2337 -280
rect 2403 -246 2495 -240
rect 2403 -280 2415 -246
rect 2483 -280 2495 -246
rect 2403 -286 2495 -280
rect 2561 -246 2653 -240
rect 2561 -280 2573 -246
rect 2641 -280 2653 -246
rect 2561 -286 2653 -280
rect 2719 -246 2811 -240
rect 2719 -280 2731 -246
rect 2799 -280 2811 -246
rect 2719 -286 2811 -280
rect 2877 -246 2969 -240
rect 2877 -280 2889 -246
rect 2957 -280 2969 -246
rect 2877 -286 2969 -280
rect 3035 -246 3127 -240
rect 3035 -280 3047 -246
rect 3115 -280 3127 -246
rect 3035 -286 3127 -280
rect -3183 -330 -3137 -318
rect -3183 -506 -3177 -330
rect -3143 -506 -3137 -330
rect -3183 -518 -3137 -506
rect -3025 -330 -2979 -318
rect -3025 -506 -3019 -330
rect -2985 -506 -2979 -330
rect -3025 -518 -2979 -506
rect -2867 -330 -2821 -318
rect -2867 -506 -2861 -330
rect -2827 -506 -2821 -330
rect -2867 -518 -2821 -506
rect -2709 -330 -2663 -318
rect -2709 -506 -2703 -330
rect -2669 -506 -2663 -330
rect -2709 -518 -2663 -506
rect -2551 -330 -2505 -318
rect -2551 -506 -2545 -330
rect -2511 -506 -2505 -330
rect -2551 -518 -2505 -506
rect -2393 -330 -2347 -318
rect -2393 -506 -2387 -330
rect -2353 -506 -2347 -330
rect -2393 -518 -2347 -506
rect -2235 -330 -2189 -318
rect -2235 -506 -2229 -330
rect -2195 -506 -2189 -330
rect -2235 -518 -2189 -506
rect -2077 -330 -2031 -318
rect -2077 -506 -2071 -330
rect -2037 -506 -2031 -330
rect -2077 -518 -2031 -506
rect -1919 -330 -1873 -318
rect -1919 -506 -1913 -330
rect -1879 -506 -1873 -330
rect -1919 -518 -1873 -506
rect -1761 -330 -1715 -318
rect -1761 -506 -1755 -330
rect -1721 -506 -1715 -330
rect -1761 -518 -1715 -506
rect -1603 -330 -1557 -318
rect -1603 -506 -1597 -330
rect -1563 -506 -1557 -330
rect -1603 -518 -1557 -506
rect -1445 -330 -1399 -318
rect -1445 -506 -1439 -330
rect -1405 -506 -1399 -330
rect -1445 -518 -1399 -506
rect -1287 -330 -1241 -318
rect -1287 -506 -1281 -330
rect -1247 -506 -1241 -330
rect -1287 -518 -1241 -506
rect -1129 -330 -1083 -318
rect -1129 -506 -1123 -330
rect -1089 -506 -1083 -330
rect -1129 -518 -1083 -506
rect -971 -330 -925 -318
rect -971 -506 -965 -330
rect -931 -506 -925 -330
rect -971 -518 -925 -506
rect -813 -330 -767 -318
rect -813 -506 -807 -330
rect -773 -506 -767 -330
rect -813 -518 -767 -506
rect -655 -330 -609 -318
rect -655 -506 -649 -330
rect -615 -506 -609 -330
rect -655 -518 -609 -506
rect -497 -330 -451 -318
rect -497 -506 -491 -330
rect -457 -506 -451 -330
rect -497 -518 -451 -506
rect -339 -330 -293 -318
rect -339 -506 -333 -330
rect -299 -506 -293 -330
rect -339 -518 -293 -506
rect -181 -330 -135 -318
rect -181 -506 -175 -330
rect -141 -506 -135 -330
rect -181 -518 -135 -506
rect -23 -330 23 -318
rect -23 -506 -17 -330
rect 17 -506 23 -330
rect -23 -518 23 -506
rect 135 -330 181 -318
rect 135 -506 141 -330
rect 175 -506 181 -330
rect 135 -518 181 -506
rect 293 -330 339 -318
rect 293 -506 299 -330
rect 333 -506 339 -330
rect 293 -518 339 -506
rect 451 -330 497 -318
rect 451 -506 457 -330
rect 491 -506 497 -330
rect 451 -518 497 -506
rect 609 -330 655 -318
rect 609 -506 615 -330
rect 649 -506 655 -330
rect 609 -518 655 -506
rect 767 -330 813 -318
rect 767 -506 773 -330
rect 807 -506 813 -330
rect 767 -518 813 -506
rect 925 -330 971 -318
rect 925 -506 931 -330
rect 965 -506 971 -330
rect 925 -518 971 -506
rect 1083 -330 1129 -318
rect 1083 -506 1089 -330
rect 1123 -506 1129 -330
rect 1083 -518 1129 -506
rect 1241 -330 1287 -318
rect 1241 -506 1247 -330
rect 1281 -506 1287 -330
rect 1241 -518 1287 -506
rect 1399 -330 1445 -318
rect 1399 -506 1405 -330
rect 1439 -506 1445 -330
rect 1399 -518 1445 -506
rect 1557 -330 1603 -318
rect 1557 -506 1563 -330
rect 1597 -506 1603 -330
rect 1557 -518 1603 -506
rect 1715 -330 1761 -318
rect 1715 -506 1721 -330
rect 1755 -506 1761 -330
rect 1715 -518 1761 -506
rect 1873 -330 1919 -318
rect 1873 -506 1879 -330
rect 1913 -506 1919 -330
rect 1873 -518 1919 -506
rect 2031 -330 2077 -318
rect 2031 -506 2037 -330
rect 2071 -506 2077 -330
rect 2031 -518 2077 -506
rect 2189 -330 2235 -318
rect 2189 -506 2195 -330
rect 2229 -506 2235 -330
rect 2189 -518 2235 -506
rect 2347 -330 2393 -318
rect 2347 -506 2353 -330
rect 2387 -506 2393 -330
rect 2347 -518 2393 -506
rect 2505 -330 2551 -318
rect 2505 -506 2511 -330
rect 2545 -506 2551 -330
rect 2505 -518 2551 -506
rect 2663 -330 2709 -318
rect 2663 -506 2669 -330
rect 2703 -506 2709 -330
rect 2663 -518 2709 -506
rect 2821 -330 2867 -318
rect 2821 -506 2827 -330
rect 2861 -506 2867 -330
rect 2821 -518 2867 -506
rect 2979 -330 3025 -318
rect 2979 -506 2985 -330
rect 3019 -506 3025 -330
rect 2979 -518 3025 -506
rect 3137 -330 3183 -318
rect 3137 -506 3143 -330
rect 3177 -506 3183 -330
rect 3137 -518 3183 -506
rect -3127 -556 -3035 -550
rect -3127 -590 -3115 -556
rect -3047 -590 -3035 -556
rect -3127 -596 -3035 -590
rect -2969 -556 -2877 -550
rect -2969 -590 -2957 -556
rect -2889 -590 -2877 -556
rect -2969 -596 -2877 -590
rect -2811 -556 -2719 -550
rect -2811 -590 -2799 -556
rect -2731 -590 -2719 -556
rect -2811 -596 -2719 -590
rect -2653 -556 -2561 -550
rect -2653 -590 -2641 -556
rect -2573 -590 -2561 -556
rect -2653 -596 -2561 -590
rect -2495 -556 -2403 -550
rect -2495 -590 -2483 -556
rect -2415 -590 -2403 -556
rect -2495 -596 -2403 -590
rect -2337 -556 -2245 -550
rect -2337 -590 -2325 -556
rect -2257 -590 -2245 -556
rect -2337 -596 -2245 -590
rect -2179 -556 -2087 -550
rect -2179 -590 -2167 -556
rect -2099 -590 -2087 -556
rect -2179 -596 -2087 -590
rect -2021 -556 -1929 -550
rect -2021 -590 -2009 -556
rect -1941 -590 -1929 -556
rect -2021 -596 -1929 -590
rect -1863 -556 -1771 -550
rect -1863 -590 -1851 -556
rect -1783 -590 -1771 -556
rect -1863 -596 -1771 -590
rect -1705 -556 -1613 -550
rect -1705 -590 -1693 -556
rect -1625 -590 -1613 -556
rect -1705 -596 -1613 -590
rect -1547 -556 -1455 -550
rect -1547 -590 -1535 -556
rect -1467 -590 -1455 -556
rect -1547 -596 -1455 -590
rect -1389 -556 -1297 -550
rect -1389 -590 -1377 -556
rect -1309 -590 -1297 -556
rect -1389 -596 -1297 -590
rect -1231 -556 -1139 -550
rect -1231 -590 -1219 -556
rect -1151 -590 -1139 -556
rect -1231 -596 -1139 -590
rect -1073 -556 -981 -550
rect -1073 -590 -1061 -556
rect -993 -590 -981 -556
rect -1073 -596 -981 -590
rect -915 -556 -823 -550
rect -915 -590 -903 -556
rect -835 -590 -823 -556
rect -915 -596 -823 -590
rect -757 -556 -665 -550
rect -757 -590 -745 -556
rect -677 -590 -665 -556
rect -757 -596 -665 -590
rect -599 -556 -507 -550
rect -599 -590 -587 -556
rect -519 -590 -507 -556
rect -599 -596 -507 -590
rect -441 -556 -349 -550
rect -441 -590 -429 -556
rect -361 -590 -349 -556
rect -441 -596 -349 -590
rect -283 -556 -191 -550
rect -283 -590 -271 -556
rect -203 -590 -191 -556
rect -283 -596 -191 -590
rect -125 -556 -33 -550
rect -125 -590 -113 -556
rect -45 -590 -33 -556
rect -125 -596 -33 -590
rect 33 -556 125 -550
rect 33 -590 45 -556
rect 113 -590 125 -556
rect 33 -596 125 -590
rect 191 -556 283 -550
rect 191 -590 203 -556
rect 271 -590 283 -556
rect 191 -596 283 -590
rect 349 -556 441 -550
rect 349 -590 361 -556
rect 429 -590 441 -556
rect 349 -596 441 -590
rect 507 -556 599 -550
rect 507 -590 519 -556
rect 587 -590 599 -556
rect 507 -596 599 -590
rect 665 -556 757 -550
rect 665 -590 677 -556
rect 745 -590 757 -556
rect 665 -596 757 -590
rect 823 -556 915 -550
rect 823 -590 835 -556
rect 903 -590 915 -556
rect 823 -596 915 -590
rect 981 -556 1073 -550
rect 981 -590 993 -556
rect 1061 -590 1073 -556
rect 981 -596 1073 -590
rect 1139 -556 1231 -550
rect 1139 -590 1151 -556
rect 1219 -590 1231 -556
rect 1139 -596 1231 -590
rect 1297 -556 1389 -550
rect 1297 -590 1309 -556
rect 1377 -590 1389 -556
rect 1297 -596 1389 -590
rect 1455 -556 1547 -550
rect 1455 -590 1467 -556
rect 1535 -590 1547 -556
rect 1455 -596 1547 -590
rect 1613 -556 1705 -550
rect 1613 -590 1625 -556
rect 1693 -590 1705 -556
rect 1613 -596 1705 -590
rect 1771 -556 1863 -550
rect 1771 -590 1783 -556
rect 1851 -590 1863 -556
rect 1771 -596 1863 -590
rect 1929 -556 2021 -550
rect 1929 -590 1941 -556
rect 2009 -590 2021 -556
rect 1929 -596 2021 -590
rect 2087 -556 2179 -550
rect 2087 -590 2099 -556
rect 2167 -590 2179 -556
rect 2087 -596 2179 -590
rect 2245 -556 2337 -550
rect 2245 -590 2257 -556
rect 2325 -590 2337 -556
rect 2245 -596 2337 -590
rect 2403 -556 2495 -550
rect 2403 -590 2415 -556
rect 2483 -590 2495 -556
rect 2403 -596 2495 -590
rect 2561 -556 2653 -550
rect 2561 -590 2573 -556
rect 2641 -590 2653 -556
rect 2561 -596 2653 -590
rect 2719 -556 2811 -550
rect 2719 -590 2731 -556
rect 2799 -590 2811 -556
rect 2719 -596 2811 -590
rect 2877 -556 2969 -550
rect 2877 -590 2889 -556
rect 2957 -590 2969 -556
rect 2877 -596 2969 -590
rect 3035 -556 3127 -550
rect 3035 -590 3047 -556
rect 3115 -590 3127 -556
rect 3035 -596 3127 -590
<< properties >>
string FIXED_BBOX -3294 -711 3294 711
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 3 nf 40 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
